
module DPA_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4;
  wire   [19:1] carry;

  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  CLKBUFX3 U1 ( .A(B[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[1]), .B(A[1]), .Y(n1) );
  NAND2X1 U3 ( .A(B[18]), .B(n2), .Y(n4) );
  AND2X2 U4 ( .A(B[17]), .B(carry[17]), .Y(n2) );
  XOR2XL U5 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  XNOR2X1 U6 ( .A(B[19]), .B(n4), .Y(SUM[19]) );
  XOR2X1 U7 ( .A(B[18]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U8 ( .A(B[17]), .B(carry[17]), .Y(SUM[17]) );
endmodule


module DPA_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [19:1] carry;

  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  CLKBUFX3 U1 ( .A(B[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U3 ( .A(B[19]), .B(n2), .Y(SUM[19]) );
  AND2X2 U4 ( .A(B[18]), .B(n3), .Y(n2) );
  AND2X2 U5 ( .A(B[17]), .B(carry[17]), .Y(n3) );
  XOR2XL U6 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  XOR2XL U7 ( .A(B[18]), .B(n3), .Y(SUM[18]) );
  XOR2XL U8 ( .A(B[17]), .B(carry[17]), .Y(SUM[17]) );
endmodule


module DPA_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_inc_2 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_inc_3 ( A, SUM );
  input [19:0] A;
  output [19:0] SUM;

  wire   [19:2] carry;

  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  XOR2X1 U1 ( .A(carry[19]), .B(A[19]), .Y(SUM[19]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_3 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2XL U2 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  AND2X2 U3 ( .A(B[18]), .B(carry[18]), .Y(n2) );
  XOR2X1 U4 ( .A(B[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKBUFX3 U5 ( .A(B[0]), .Y(SUM[0]) );
  XOR2X1 U6 ( .A(B[19]), .B(n2), .Y(SUM[19]) );
  CLKBUFX2 U7 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module DPA_DW01_add_4 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [15:1] carry;
  assign carry[2] = A[1];

  AND2X2 U1 ( .A(A[2]), .B(carry[2]), .Y(n1) );
  AND2X2 U2 ( .A(A[3]), .B(n1), .Y(n2) );
  AND2X2 U3 ( .A(A[4]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[5]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[6]), .B(n4), .Y(n5) );
  OR2X1 U6 ( .A(A[7]), .B(n5), .Y(carry[8]) );
  AND2X2 U7 ( .A(A[8]), .B(carry[8]), .Y(n6) );
  AND2X2 U8 ( .A(A[9]), .B(n6), .Y(n7) );
  AND2X2 U9 ( .A(A[10]), .B(n7), .Y(n8) );
  AND2X2 U10 ( .A(A[11]), .B(n8), .Y(n9) );
  AND2X2 U11 ( .A(A[12]), .B(n9), .Y(n10) );
  AND2X2 U12 ( .A(A[13]), .B(n10), .Y(n11) );
  AND2X2 U13 ( .A(A[14]), .B(n11), .Y(n12) );
  XOR2XL U14 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  XOR2XL U15 ( .A(A[3]), .B(n1), .Y(SUM[3]) );
  XOR2XL U16 ( .A(A[4]), .B(n2), .Y(SUM[4]) );
  XOR2XL U17 ( .A(A[5]), .B(n3), .Y(SUM[5]) );
  XOR2XL U18 ( .A(A[6]), .B(n4), .Y(SUM[6]) );
  XNOR2XL U19 ( .A(A[7]), .B(n5), .Y(SUM[7]) );
  XOR2XL U20 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U21 ( .A(A[9]), .B(n6), .Y(SUM[9]) );
  XOR2XL U22 ( .A(A[10]), .B(n7), .Y(SUM[10]) );
  XOR2XL U23 ( .A(A[11]), .B(n8), .Y(SUM[11]) );
  XOR2XL U24 ( .A(A[12]), .B(n9), .Y(SUM[12]) );
  XOR2XL U25 ( .A(A[13]), .B(n10), .Y(SUM[13]) );
  XOR2XL U26 ( .A(A[14]), .B(n11), .Y(SUM[14]) );
  INVXL U27 ( .A(carry[2]), .Y(SUM[1]) );
  XOR2XL U28 ( .A(A[15]), .B(n12), .Y(SUM[15]) );
  CLKBUFX2 U29 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_5 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   \carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14;
  assign \carry[2]  = A[1];

  AND2X2 U1 ( .A(A[2]), .B(\carry[2] ), .Y(n1) );
  AND2X2 U2 ( .A(A[4]), .B(n12), .Y(n2) );
  AND2X2 U3 ( .A(A[5]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[6]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[7]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[8]), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(A[10]), .B(n11), .Y(n7) );
  AND2X2 U8 ( .A(A[11]), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(A[12]), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(A[13]), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(A[9]), .B(n6), .Y(n11) );
  XOR2X1 U12 ( .A(A[3]), .B(n1), .Y(SUM[3]) );
  AND2X2 U13 ( .A(A[3]), .B(n1), .Y(n12) );
  XOR2X1 U14 ( .A(A[5]), .B(n2), .Y(SUM[5]) );
  XOR2X1 U15 ( .A(A[6]), .B(n3), .Y(SUM[6]) );
  XOR2X1 U16 ( .A(A[7]), .B(n4), .Y(SUM[7]) );
  XOR2X1 U17 ( .A(A[8]), .B(n5), .Y(SUM[8]) );
  XOR2X1 U18 ( .A(A[9]), .B(n6), .Y(SUM[9]) );
  XOR2X1 U19 ( .A(A[11]), .B(n7), .Y(SUM[11]) );
  XOR2X1 U20 ( .A(A[12]), .B(n8), .Y(SUM[12]) );
  XOR2X1 U21 ( .A(A[13]), .B(n9), .Y(SUM[13]) );
  XOR2X1 U22 ( .A(A[14]), .B(n10), .Y(SUM[14]) );
  XNOR2X1 U23 ( .A(A[15]), .B(n14), .Y(SUM[15]) );
  NAND2X1 U24 ( .A(A[14]), .B(n10), .Y(n14) );
  XOR2X1 U25 ( .A(A[10]), .B(n11), .Y(SUM[10]) );
  INVX1 U26 ( .A(\carry[2] ), .Y(SUM[1]) );
  XOR2XL U27 ( .A(A[2]), .B(\carry[2] ), .Y(SUM[2]) );
  XOR2X1 U28 ( .A(A[4]), .B(n12), .Y(SUM[4]) );
  CLKBUFX2 U29 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_6 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [24:1] carry;

  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module DPA_DW01_add_7 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U2 ( .A(B[18]), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(B[17]), .B(carry[17]), .Y(n3) );
  XOR2XL U4 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U5 ( .A(B[0]), .Y(SUM[0]) );
  XOR2X1 U6 ( .A(B[19]), .B(n2), .Y(SUM[19]) );
  XOR2X1 U7 ( .A(B[18]), .B(n3), .Y(SUM[18]) );
  XOR2X1 U8 ( .A(B[17]), .B(carry[17]), .Y(SUM[17]) );
endmodule


module DPA_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [16:0] carry;
  assign carry[1] = A[0];

  AND2X2 U1 ( .A(A[1]), .B(carry[1]), .Y(n1) );
  AND2X2 U2 ( .A(A[2]), .B(n1), .Y(n2) );
  AND2X2 U3 ( .A(A[3]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[4]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[5]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[6]), .B(n5), .Y(n6) );
  OR2X1 U7 ( .A(A[7]), .B(n6), .Y(carry[8]) );
  OR2X1 U8 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  OR2X1 U9 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
  OR2X1 U10 ( .A(A[11]), .B(carry[11]), .Y(carry[12]) );
  OR2X1 U11 ( .A(A[12]), .B(carry[12]), .Y(carry[13]) );
  OR2X1 U12 ( .A(A[13]), .B(carry[13]), .Y(carry[14]) );
  OR2X1 U13 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  XOR2XL U14 ( .A(A[1]), .B(carry[1]), .Y(DIFF[1]) );
  XOR2X1 U15 ( .A(A[2]), .B(n1), .Y(DIFF[2]) );
  XOR2X1 U16 ( .A(A[3]), .B(n2), .Y(DIFF[3]) );
  XOR2X1 U17 ( .A(A[4]), .B(n3), .Y(DIFF[4]) );
  XOR2X1 U18 ( .A(A[5]), .B(n4), .Y(DIFF[5]) );
  XOR2X1 U19 ( .A(A[6]), .B(n5), .Y(DIFF[6]) );
  XNOR2X1 U20 ( .A(A[7]), .B(n6), .Y(DIFF[7]) );
  XNOR2X1 U21 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2X1 U22 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2X1 U23 ( .A(A[11]), .B(carry[11]), .Y(DIFF[11]) );
  XNOR2X1 U24 ( .A(A[12]), .B(carry[12]), .Y(DIFF[12]) );
  XNOR2X1 U25 ( .A(A[13]), .B(carry[13]), .Y(DIFF[13]) );
  XNOR2X1 U26 ( .A(A[14]), .B(carry[14]), .Y(DIFF[14]) );
  XNOR2X1 U27 ( .A(A[15]), .B(carry[15]), .Y(DIFF[15]) );
  NAND2X1 U28 ( .A(n7), .B(n8), .Y(carry[15]) );
  INVX1 U29 ( .A(A[14]), .Y(n7) );
  CLKINVX1 U30 ( .A(carry[14]), .Y(n8) );
  XNOR2X1 U31 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  CLKINVX1 U32 ( .A(carry[1]), .Y(DIFF[0]) );
endmodule


module DPA_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [20:0] carry;
  wire   [19:0] B_not;

  ADDFXL U2_4 ( .A(A[4]), .B(B_not[4]), .CI(carry[4]), .CO(carry[5]), .S(
        DIFF[4]) );
  ADDFXL U2_5 ( .A(A[5]), .B(B_not[5]), .CI(carry[5]), .CO(carry[6]), .S(
        DIFF[5]) );
  ADDFXL U2_6 ( .A(A[6]), .B(B_not[6]), .CI(carry[6]), .CO(carry[7]), .S(
        DIFF[6]) );
  ADDFXL U2_7 ( .A(A[7]), .B(B_not[7]), .CI(carry[7]), .CO(carry[8]), .S(
        DIFF[7]) );
  ADDFXL U2_8 ( .A(A[8]), .B(B_not[8]), .CI(carry[8]), .CO(carry[9]), .S(
        DIFF[8]) );
  ADDFXL U2_9 ( .A(A[9]), .B(B_not[9]), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  ADDFXL U2_2 ( .A(A[2]), .B(B_not[2]), .CI(carry[2]), .CO(carry[3]), .S(
        DIFF[2]) );
  ADDFXL U2_1 ( .A(A[1]), .B(B_not[1]), .CI(carry[1]), .CO(carry[2]), .S(
        DIFF[1]) );
  ADDFXL U2_3 ( .A(A[3]), .B(B_not[3]), .CI(carry[3]), .CO(carry[4]), .S(
        DIFF[3]) );
  INVXL U1 ( .A(A[0]), .Y(n3) );
  OR2X1 U2 ( .A(A[17]), .B(carry[17]), .Y(carry[18]) );
  OR2X1 U3 ( .A(A[16]), .B(carry[16]), .Y(carry[17]) );
  OR2X1 U4 ( .A(A[15]), .B(carry[15]), .Y(carry[16]) );
  OR2X1 U5 ( .A(A[14]), .B(carry[14]), .Y(carry[15]) );
  OR2X1 U6 ( .A(A[13]), .B(carry[13]), .Y(carry[14]) );
  OR2X1 U7 ( .A(A[12]), .B(carry[12]), .Y(carry[13]) );
  OR2X1 U8 ( .A(A[11]), .B(carry[11]), .Y(carry[12]) );
  OR2X1 U9 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
  NAND2X1 U10 ( .A(B[0]), .B(n3), .Y(carry[1]) );
  XNOR2X1 U11 ( .A(A[19]), .B(carry[19]), .Y(DIFF[19]) );
  NAND2X1 U12 ( .A(n1), .B(n2), .Y(carry[19]) );
  CLKINVX1 U13 ( .A(A[18]), .Y(n1) );
  CLKINVX1 U14 ( .A(carry[18]), .Y(n2) );
  XNOR2X1 U15 ( .A(A[18]), .B(carry[18]), .Y(DIFF[18]) );
  XNOR2X1 U16 ( .A(A[17]), .B(carry[17]), .Y(DIFF[17]) );
  XNOR2X1 U17 ( .A(A[16]), .B(carry[16]), .Y(DIFF[16]) );
  XNOR2XL U18 ( .A(A[15]), .B(carry[15]), .Y(DIFF[15]) );
  XNOR2XL U19 ( .A(A[14]), .B(carry[14]), .Y(DIFF[14]) );
  XNOR2XL U20 ( .A(A[13]), .B(carry[13]), .Y(DIFF[13]) );
  XNOR2X1 U21 ( .A(A[12]), .B(carry[12]), .Y(DIFF[12]) );
  XNOR2X1 U22 ( .A(A[11]), .B(carry[11]), .Y(DIFF[11]) );
  XNOR2X1 U23 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  XNOR2XL U24 ( .A(B_not[0]), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U25 ( .A(B[9]), .Y(B_not[9]) );
  CLKINVX1 U26 ( .A(B[8]), .Y(B_not[8]) );
  CLKINVX1 U27 ( .A(B[7]), .Y(B_not[7]) );
  CLKINVX1 U28 ( .A(B[6]), .Y(B_not[6]) );
  CLKINVX1 U29 ( .A(B[5]), .Y(B_not[5]) );
  CLKINVX1 U30 ( .A(B[4]), .Y(B_not[4]) );
  CLKINVX1 U31 ( .A(B[3]), .Y(B_not[3]) );
  CLKINVX1 U32 ( .A(B[2]), .Y(B_not[2]) );
  CLKINVX1 U33 ( .A(B[1]), .Y(B_not[1]) );
  CLKINVX1 U34 ( .A(B[0]), .Y(B_not[0]) );
endmodule


module DPA_DW01_add_14 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [20:1] carry;
  assign carry[1] = A[0];

  OR2X1 U1 ( .A(A[4]), .B(carry[4]), .Y(carry[5]) );
  OR2X1 U2 ( .A(A[15]), .B(carry[15]), .Y(carry[16]) );
  OR2X1 U3 ( .A(A[14]), .B(carry[14]), .Y(carry[15]) );
  OR2X1 U4 ( .A(A[1]), .B(carry[1]), .Y(carry[2]) );
  OR2X1 U5 ( .A(A[12]), .B(carry[12]), .Y(carry[13]) );
  OR2X1 U6 ( .A(A[11]), .B(carry[11]), .Y(carry[12]) );
  OR2X1 U7 ( .A(A[2]), .B(carry[2]), .Y(carry[3]) );
  OR2X1 U8 ( .A(A[13]), .B(carry[13]), .Y(carry[14]) );
  OR2X1 U9 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
  OR2X1 U10 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  OR2X1 U11 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  OR2X1 U12 ( .A(A[7]), .B(carry[7]), .Y(carry[8]) );
  OR2X1 U13 ( .A(A[6]), .B(carry[6]), .Y(carry[7]) );
  OR2X1 U14 ( .A(A[5]), .B(carry[5]), .Y(carry[6]) );
  OR2X1 U15 ( .A(A[3]), .B(carry[3]), .Y(carry[4]) );
  AND2X2 U16 ( .A(A[17]), .B(n3), .Y(n1) );
  XOR2X1 U17 ( .A(A[16]), .B(carry[16]), .Y(SUM[16]) );
  XNOR2X1 U18 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  AND2X2 U19 ( .A(A[18]), .B(n1), .Y(n2) );
  AND2X2 U20 ( .A(A[16]), .B(carry[16]), .Y(n3) );
  XOR2X1 U21 ( .A(A[19]), .B(n2), .Y(SUM[19]) );
  XNOR2X1 U22 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  XNOR2X1 U23 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  XNOR2X1 U24 ( .A(A[13]), .B(carry[13]), .Y(SUM[13]) );
  XNOR2X1 U25 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XNOR2X1 U26 ( .A(A[3]), .B(carry[3]), .Y(SUM[3]) );
  XNOR2X1 U27 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XNOR2X1 U28 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  XNOR2X1 U29 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  XNOR2X1 U30 ( .A(A[9]), .B(carry[9]), .Y(SUM[9]) );
  XNOR2X1 U31 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XNOR2X1 U32 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  XNOR2X1 U33 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XNOR2X1 U34 ( .A(A[1]), .B(carry[1]), .Y(SUM[1]) );
  XNOR2X1 U35 ( .A(A[4]), .B(carry[4]), .Y(SUM[4]) );
  XOR2X1 U36 ( .A(A[18]), .B(n1), .Y(SUM[18]) );
  AND2X2 U37 ( .A(A[19]), .B(n2), .Y(SUM[20]) );
  XOR2X1 U38 ( .A(A[17]), .B(n3), .Y(SUM[17]) );
  CLKINVX1 U39 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_15 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(A[18]), .B(n13), .Y(SUM[18]) );
  AND2X2 U2 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U3 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  XOR2X1 U4 ( .A(A[17]), .B(n14), .Y(SUM[17]) );
  AND2X2 U5 ( .A(A[6]), .B(n3), .Y(n2) );
  AND2X2 U6 ( .A(A[5]), .B(carry[5]), .Y(n3) );
  AND2X2 U7 ( .A(A[15]), .B(n5), .Y(n4) );
  AND2X2 U8 ( .A(A[14]), .B(n6), .Y(n5) );
  AND2X2 U9 ( .A(A[13]), .B(n7), .Y(n6) );
  AND2X2 U10 ( .A(A[12]), .B(n8), .Y(n7) );
  AND2X2 U11 ( .A(A[11]), .B(n9), .Y(n8) );
  AND2X2 U12 ( .A(A[10]), .B(n10), .Y(n9) );
  AND2X2 U13 ( .A(A[9]), .B(n11), .Y(n10) );
  AND2X2 U14 ( .A(A[8]), .B(n12), .Y(n11) );
  AND2X2 U15 ( .A(A[7]), .B(n2), .Y(n12) );
  XOR2X1 U16 ( .A(A[7]), .B(n2), .Y(SUM[7]) );
  XOR2X1 U17 ( .A(A[6]), .B(n3), .Y(SUM[6]) );
  XOR2X1 U18 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  AND2X2 U19 ( .A(A[17]), .B(n14), .Y(n13) );
  AND2X2 U20 ( .A(A[16]), .B(n4), .Y(n14) );
  XOR2X1 U21 ( .A(A[16]), .B(n4), .Y(SUM[16]) );
  XOR2X1 U22 ( .A(A[15]), .B(n5), .Y(SUM[15]) );
  XOR2X1 U23 ( .A(A[14]), .B(n6), .Y(SUM[14]) );
  XOR2X1 U24 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U25 ( .A(A[12]), .B(n8), .Y(SUM[12]) );
  XOR2X1 U26 ( .A(A[11]), .B(n9), .Y(SUM[11]) );
  XOR2X1 U27 ( .A(A[10]), .B(n10), .Y(SUM[10]) );
  XOR2X1 U28 ( .A(A[9]), .B(n11), .Y(SUM[9]) );
  XOR2X1 U29 ( .A(A[8]), .B(n12), .Y(SUM[8]) );
  CLKBUFX2 U30 ( .A(A[0]), .Y(SUM[0]) );
  XNOR2X1 U31 ( .A(A[19]), .B(n16), .Y(SUM[19]) );
  NAND2X1 U32 ( .A(A[18]), .B(n13), .Y(n16) );
endmodule


module DPA_DW01_add_16 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [19:1] carry;
  assign carry[1] = B[0];

  XOR2X1 U1 ( .A(B[18]), .B(n14), .Y(SUM[18]) );
  XOR2X1 U2 ( .A(B[17]), .B(n15), .Y(SUM[17]) );
  AND2X2 U3 ( .A(B[1]), .B(carry[1]), .Y(n1) );
  AND2X2 U4 ( .A(B[6]), .B(n3), .Y(n2) );
  AND2X2 U5 ( .A(B[5]), .B(n4), .Y(n3) );
  AND2X2 U6 ( .A(B[4]), .B(n5), .Y(n4) );
  AND2X2 U7 ( .A(B[3]), .B(n6), .Y(n5) );
  AND2X2 U8 ( .A(B[2]), .B(n1), .Y(n6) );
  XOR2X1 U9 ( .A(B[2]), .B(n1), .Y(SUM[2]) );
  AND2X2 U10 ( .A(B[15]), .B(n8), .Y(n7) );
  AND2X2 U11 ( .A(B[14]), .B(n9), .Y(n8) );
  AND2X2 U12 ( .A(B[13]), .B(n10), .Y(n9) );
  AND2X2 U13 ( .A(B[12]), .B(n11), .Y(n10) );
  AND2X2 U14 ( .A(B[11]), .B(n12), .Y(n11) );
  AND2X2 U15 ( .A(B[10]), .B(carry[10]), .Y(n12) );
  OR2X1 U16 ( .A(B[9]), .B(carry[9]), .Y(carry[10]) );
  OR2X1 U17 ( .A(B[8]), .B(n13), .Y(carry[9]) );
  AND2X2 U18 ( .A(B[7]), .B(n2), .Y(n13) );
  XOR2X1 U19 ( .A(B[7]), .B(n2), .Y(SUM[7]) );
  XOR2X1 U20 ( .A(B[6]), .B(n3), .Y(SUM[6]) );
  XOR2X1 U21 ( .A(B[5]), .B(n4), .Y(SUM[5]) );
  XOR2X1 U22 ( .A(B[4]), .B(n5), .Y(SUM[4]) );
  XOR2X1 U23 ( .A(B[3]), .B(n6), .Y(SUM[3]) );
  AND2X2 U24 ( .A(B[17]), .B(n15), .Y(n14) );
  AND2X2 U25 ( .A(B[16]), .B(n7), .Y(n15) );
  XOR2X1 U26 ( .A(B[16]), .B(n7), .Y(SUM[16]) );
  XOR2X1 U27 ( .A(B[15]), .B(n8), .Y(SUM[15]) );
  XOR2X1 U28 ( .A(B[14]), .B(n9), .Y(SUM[14]) );
  XOR2X1 U29 ( .A(B[13]), .B(n10), .Y(SUM[13]) );
  XOR2X1 U30 ( .A(B[12]), .B(n11), .Y(SUM[12]) );
  XOR2X1 U31 ( .A(B[11]), .B(n12), .Y(SUM[11]) );
  XOR2X1 U32 ( .A(B[10]), .B(carry[10]), .Y(SUM[10]) );
  XNOR2X1 U33 ( .A(B[9]), .B(carry[9]), .Y(SUM[9]) );
  XNOR2X1 U34 ( .A(B[8]), .B(n13), .Y(SUM[8]) );
  XOR2X1 U35 ( .A(B[1]), .B(carry[1]), .Y(SUM[1]) );
  XNOR2X1 U36 ( .A(B[19]), .B(n16), .Y(SUM[19]) );
  NAND2X1 U37 ( .A(B[18]), .B(n14), .Y(n16) );
  CLKINVX1 U38 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_17 ( A, B, CI, SUM, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [25:1] carry;

  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_18 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [19:1] carry;
  assign carry[1] = B[0];

  XOR2X1 U1 ( .A(B[9]), .B(carry[9]), .Y(SUM[9]) );
  XOR2X1 U2 ( .A(B[1]), .B(carry[1]), .Y(SUM[1]) );
  XOR2X1 U3 ( .A(B[12]), .B(n11), .Y(SUM[12]) );
  XOR2X1 U4 ( .A(B[7]), .B(n2), .Y(SUM[7]) );
  XOR2X1 U5 ( .A(B[6]), .B(n3), .Y(SUM[6]) );
  XOR2X1 U6 ( .A(B[5]), .B(n4), .Y(SUM[5]) );
  XOR2X1 U7 ( .A(B[15]), .B(n8), .Y(SUM[15]) );
  XOR2X1 U8 ( .A(B[14]), .B(n9), .Y(SUM[14]) );
  XOR2X1 U9 ( .A(B[13]), .B(n10), .Y(SUM[13]) );
  XOR2X1 U10 ( .A(B[11]), .B(n12), .Y(SUM[11]) );
  XOR2X1 U11 ( .A(B[10]), .B(n13), .Y(SUM[10]) );
  XOR2X1 U12 ( .A(B[16]), .B(n7), .Y(SUM[16]) );
  XNOR2X1 U13 ( .A(B[8]), .B(n14), .Y(SUM[8]) );
  XOR2X1 U14 ( .A(B[17]), .B(n16), .Y(SUM[17]) );
  AND2X2 U15 ( .A(B[1]), .B(carry[1]), .Y(n1) );
  AND2X2 U16 ( .A(B[6]), .B(n3), .Y(n2) );
  AND2X2 U17 ( .A(B[5]), .B(n4), .Y(n3) );
  AND2X2 U18 ( .A(B[4]), .B(n5), .Y(n4) );
  AND2X2 U19 ( .A(B[3]), .B(n6), .Y(n5) );
  AND2X2 U20 ( .A(B[2]), .B(n1), .Y(n6) );
  XOR2X1 U21 ( .A(B[2]), .B(n1), .Y(SUM[2]) );
  AND2X2 U22 ( .A(B[15]), .B(n8), .Y(n7) );
  AND2X2 U23 ( .A(B[14]), .B(n9), .Y(n8) );
  AND2X2 U24 ( .A(B[13]), .B(n10), .Y(n9) );
  AND2X2 U25 ( .A(B[12]), .B(n11), .Y(n10) );
  AND2X2 U26 ( .A(B[11]), .B(n12), .Y(n11) );
  AND2X2 U27 ( .A(B[10]), .B(n13), .Y(n12) );
  AND2X2 U28 ( .A(B[9]), .B(carry[9]), .Y(n13) );
  OR2X1 U29 ( .A(B[8]), .B(n14), .Y(carry[9]) );
  AND2X2 U30 ( .A(B[7]), .B(n2), .Y(n14) );
  XOR2X1 U31 ( .A(B[4]), .B(n5), .Y(SUM[4]) );
  XOR2X1 U32 ( .A(B[3]), .B(n6), .Y(SUM[3]) );
  AND2X2 U33 ( .A(B[17]), .B(n16), .Y(n15) );
  AND2X2 U34 ( .A(B[16]), .B(n7), .Y(n16) );
  XNOR2X1 U35 ( .A(B[19]), .B(n17), .Y(SUM[19]) );
  NAND2X1 U36 ( .A(B[18]), .B(n15), .Y(n17) );
  CLKXOR2X2 U37 ( .A(B[18]), .B(n15), .Y(SUM[18]) );
  CLKINVX1 U38 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_19 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [15:1] carry;
  assign carry[1] = A[0];

  AND2X2 U1 ( .A(A[1]), .B(carry[1]), .Y(n1) );
  AND2X2 U2 ( .A(A[2]), .B(n1), .Y(n2) );
  AND2X2 U3 ( .A(A[3]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[4]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[5]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[6]), .B(n5), .Y(n6) );
  OR2X1 U7 ( .A(A[7]), .B(n6), .Y(carry[8]) );
  AND2X2 U8 ( .A(A[8]), .B(carry[8]), .Y(n7) );
  AND2X2 U9 ( .A(A[10]), .B(n12), .Y(n8) );
  AND2X2 U10 ( .A(A[11]), .B(n8), .Y(n9) );
  AND2X2 U11 ( .A(A[12]), .B(n9), .Y(n10) );
  AND2X2 U12 ( .A(A[13]), .B(n10), .Y(n11) );
  AND2X2 U13 ( .A(A[9]), .B(n7), .Y(n12) );
  XOR2XL U14 ( .A(A[1]), .B(carry[1]), .Y(SUM[1]) );
  XOR2X1 U15 ( .A(A[2]), .B(n1), .Y(SUM[2]) );
  XOR2X1 U16 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  XOR2X1 U17 ( .A(A[4]), .B(n3), .Y(SUM[4]) );
  XOR2X1 U18 ( .A(A[5]), .B(n4), .Y(SUM[5]) );
  XOR2X1 U19 ( .A(A[6]), .B(n5), .Y(SUM[6]) );
  XNOR2X1 U20 ( .A(A[7]), .B(n6), .Y(SUM[7]) );
  XOR2X1 U21 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U22 ( .A(A[9]), .B(n7), .Y(SUM[9]) );
  XOR2X1 U23 ( .A(A[11]), .B(n8), .Y(SUM[11]) );
  XOR2X1 U24 ( .A(A[12]), .B(n9), .Y(SUM[12]) );
  XOR2X1 U25 ( .A(A[13]), .B(n10), .Y(SUM[13]) );
  XOR2X1 U26 ( .A(A[14]), .B(n11), .Y(SUM[14]) );
  XNOR2X1 U27 ( .A(A[15]), .B(n13), .Y(SUM[15]) );
  NAND2X1 U28 ( .A(A[14]), .B(n11), .Y(n13) );
  XOR2X1 U29 ( .A(A[10]), .B(n12), .Y(SUM[10]) );
  CLKINVX1 U30 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_20 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [20:1] carry;
  assign carry[2] = A[1];

  OR2X1 U1 ( .A(A[15]), .B(carry[15]), .Y(carry[16]) );
  OR2X1 U2 ( .A(A[4]), .B(carry[4]), .Y(carry[5]) );
  OR2X1 U3 ( .A(A[3]), .B(carry[3]), .Y(carry[4]) );
  OR2X1 U4 ( .A(A[6]), .B(carry[6]), .Y(carry[7]) );
  OR2X1 U5 ( .A(A[12]), .B(carry[12]), .Y(carry[13]) );
  OR2X1 U6 ( .A(A[2]), .B(carry[2]), .Y(carry[3]) );
  OR2X1 U7 ( .A(A[14]), .B(carry[14]), .Y(carry[15]) );
  OR2X1 U8 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  OR2X1 U9 ( .A(A[7]), .B(carry[7]), .Y(carry[8]) );
  OR2X1 U10 ( .A(A[13]), .B(carry[13]), .Y(carry[14]) );
  AND2X2 U11 ( .A(A[17]), .B(n2), .Y(n1) );
  AND2X2 U12 ( .A(A[16]), .B(carry[16]), .Y(n2) );
  XOR2X1 U13 ( .A(A[16]), .B(carry[16]), .Y(SUM[16]) );
  XNOR2X1 U14 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  AND2X2 U15 ( .A(A[18]), .B(n1), .Y(n3) );
  XOR2X1 U16 ( .A(A[19]), .B(n3), .Y(SUM[19]) );
  OR2X1 U17 ( .A(A[5]), .B(carry[5]), .Y(carry[6]) );
  XNOR2X1 U18 ( .A(A[4]), .B(carry[4]), .Y(SUM[4]) );
  INVXL U19 ( .A(carry[2]), .Y(SUM[1]) );
  XNOR2X1 U20 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  XNOR2X1 U21 ( .A(A[13]), .B(carry[13]), .Y(SUM[13]) );
  XNOR2X1 U22 ( .A(A[3]), .B(carry[3]), .Y(SUM[3]) );
  OR2X1 U23 ( .A(A[11]), .B(carry[11]), .Y(carry[12]) );
  XNOR2X1 U24 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  OR2X1 U25 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
  XNOR2X1 U26 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  XNOR2X1 U27 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  OR2X1 U28 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  XNOR2X1 U29 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2X1 U30 ( .A(A[18]), .B(n1), .Y(SUM[18]) );
  XOR2X1 U31 ( .A(A[17]), .B(n2), .Y(SUM[17]) );
  AND2X2 U32 ( .A(A[19]), .B(n3), .Y(SUM[20]) );
  XNOR2X1 U33 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  CLKBUFX2 U34 ( .A(A[0]), .Y(SUM[0]) );
  XNOR2X1 U35 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XNOR2X1 U36 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  XNOR2X1 U37 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  XNOR2X1 U38 ( .A(A[9]), .B(carry[9]), .Y(SUM[9]) );
endmodule


module DPA_DW01_add_21 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [15:1] carry;
  assign carry[1] = A[0];

  AND2X2 U1 ( .A(A[1]), .B(carry[1]), .Y(n1) );
  AND2X2 U2 ( .A(A[2]), .B(n1), .Y(n2) );
  AND2X2 U3 ( .A(A[3]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[4]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[5]), .B(n4), .Y(n5) );
  OR2X1 U6 ( .A(A[6]), .B(n5), .Y(carry[7]) );
  AND2X2 U7 ( .A(A[7]), .B(carry[7]), .Y(n6) );
  AND2X2 U8 ( .A(A[8]), .B(n6), .Y(n7) );
  AND2X2 U9 ( .A(A[10]), .B(n12), .Y(n8) );
  AND2X2 U10 ( .A(A[11]), .B(n8), .Y(n9) );
  AND2X2 U11 ( .A(A[12]), .B(n9), .Y(n10) );
  AND2X2 U12 ( .A(A[13]), .B(n10), .Y(n11) );
  AND2X2 U13 ( .A(A[9]), .B(n7), .Y(n12) );
  XOR2XL U14 ( .A(A[1]), .B(carry[1]), .Y(SUM[1]) );
  XOR2X1 U15 ( .A(A[2]), .B(n1), .Y(SUM[2]) );
  XOR2X1 U16 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  XOR2X1 U17 ( .A(A[4]), .B(n3), .Y(SUM[4]) );
  XOR2X1 U18 ( .A(A[5]), .B(n4), .Y(SUM[5]) );
  XNOR2X1 U19 ( .A(A[6]), .B(n5), .Y(SUM[6]) );
  XOR2X1 U20 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  XOR2X1 U21 ( .A(A[8]), .B(n6), .Y(SUM[8]) );
  XOR2X1 U22 ( .A(A[9]), .B(n7), .Y(SUM[9]) );
  XOR2X1 U23 ( .A(A[11]), .B(n8), .Y(SUM[11]) );
  XOR2X1 U24 ( .A(A[12]), .B(n9), .Y(SUM[12]) );
  XOR2X1 U25 ( .A(A[13]), .B(n10), .Y(SUM[13]) );
  XOR2X1 U26 ( .A(A[14]), .B(n11), .Y(SUM[14]) );
  XNOR2X1 U27 ( .A(A[15]), .B(n13), .Y(SUM[15]) );
  NAND2X1 U28 ( .A(A[14]), .B(n11), .Y(n13) );
  XOR2X1 U29 ( .A(A[10]), .B(n12), .Y(SUM[10]) );
  CLKINVX1 U30 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_22 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4;
  wire   [19:1] carry;

  CMPR32X2 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .CO(carry[3]), .S(SUM[2]) );
  CMPR32X2 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CMPR32X2 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  XOR2X1 U1 ( .A(A[18]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U2 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X2 U3 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U4 ( .A(A[17]), .B(carry[17]), .Y(n2) );
  XNOR2X1 U5 ( .A(A[19]), .B(n4), .Y(SUM[19]) );
  NAND2X1 U6 ( .A(A[18]), .B(n2), .Y(n4) );
  XOR2X1 U7 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  CLKBUFX2 U8 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_inc_4 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_inc_5 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_23 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [24:1] carry;

  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module DPA_DW01_add_24 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;
  assign carry[1] = A[0];

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X1 U1 ( .A(A[18]), .B(n1), .Y(SUM[18]) );
  AND2X2 U2 ( .A(A[17]), .B(carry[17]), .Y(n1) );
  XNOR2X1 U3 ( .A(A[19]), .B(n2), .Y(SUM[19]) );
  NAND2X1 U4 ( .A(A[18]), .B(n1), .Y(n2) );
  XOR2X1 U5 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  CLKINVX1 U6 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3;
  wire   [20:0] carry;
  assign carry[2] = A[1];

  XNOR2X1 U1 ( .A(A[19]), .B(carry[19]), .Y(DIFF[19]) );
  NAND2X1 U2 ( .A(n2), .B(n3), .Y(carry[19]) );
  CLKINVX1 U3 ( .A(A[18]), .Y(n2) );
  CLKINVX1 U4 ( .A(carry[18]), .Y(n3) );
  OR2X1 U5 ( .A(A[17]), .B(carry[17]), .Y(carry[18]) );
  OR2X1 U6 ( .A(A[16]), .B(carry[16]), .Y(carry[17]) );
  OR2X1 U7 ( .A(A[15]), .B(carry[15]), .Y(carry[16]) );
  OR2X1 U8 ( .A(A[14]), .B(carry[14]), .Y(carry[15]) );
  OR2X1 U9 ( .A(A[13]), .B(carry[13]), .Y(carry[14]) );
  OR2X1 U10 ( .A(A[12]), .B(carry[12]), .Y(carry[13]) );
  OR2X1 U11 ( .A(A[11]), .B(carry[11]), .Y(carry[12]) );
  OR2X1 U12 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
  OR2X1 U13 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  OR2X1 U14 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  OR2X1 U15 ( .A(A[7]), .B(carry[7]), .Y(carry[8]) );
  OR2X1 U16 ( .A(A[6]), .B(carry[6]), .Y(carry[7]) );
  OR2X1 U17 ( .A(A[5]), .B(carry[5]), .Y(carry[6]) );
  OR2X1 U18 ( .A(A[4]), .B(carry[4]), .Y(carry[5]) );
  OR2X1 U19 ( .A(A[3]), .B(carry[3]), .Y(carry[4]) );
  OR2X1 U20 ( .A(A[2]), .B(carry[2]), .Y(carry[3]) );
  CLKBUFX3 U21 ( .A(A[0]), .Y(DIFF[0]) );
  XNOR2X1 U22 ( .A(A[2]), .B(carry[2]), .Y(DIFF[2]) );
  XNOR2X1 U23 ( .A(A[18]), .B(carry[18]), .Y(DIFF[18]) );
  XNOR2X1 U24 ( .A(A[17]), .B(carry[17]), .Y(DIFF[17]) );
  XNOR2X1 U25 ( .A(A[16]), .B(carry[16]), .Y(DIFF[16]) );
  XNOR2X1 U26 ( .A(A[15]), .B(carry[15]), .Y(DIFF[15]) );
  XNOR2X1 U27 ( .A(A[14]), .B(carry[14]), .Y(DIFF[14]) );
  XNOR2X1 U28 ( .A(A[13]), .B(carry[13]), .Y(DIFF[13]) );
  XNOR2X1 U29 ( .A(A[12]), .B(carry[12]), .Y(DIFF[12]) );
  XNOR2X1 U30 ( .A(A[11]), .B(carry[11]), .Y(DIFF[11]) );
  XNOR2X1 U31 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  XNOR2X1 U32 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2X1 U33 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2X1 U34 ( .A(A[7]), .B(carry[7]), .Y(DIFF[7]) );
  XNOR2X1 U35 ( .A(A[6]), .B(carry[6]), .Y(DIFF[6]) );
  XNOR2X1 U36 ( .A(A[5]), .B(carry[5]), .Y(DIFF[5]) );
  XNOR2X1 U37 ( .A(A[4]), .B(carry[4]), .Y(DIFF[4]) );
  XNOR2X1 U38 ( .A(A[3]), .B(carry[3]), .Y(DIFF[3]) );
  CLKINVX1 U39 ( .A(carry[2]), .Y(DIFF[1]) );
endmodule


module DPA_DW01_add_25 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n5;
  wire   [19:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  CLKINVX1 U1 ( .A(B[0]), .Y(n3) );
  AND2X2 U2 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2XL U3 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U4 ( .A(B[1]), .Y(SUM[1]) );
  CLKINVX1 U5 ( .A(n3), .Y(SUM[0]) );
  XNOR2X1 U6 ( .A(B[19]), .B(n5), .Y(SUM[19]) );
  NAND2X1 U7 ( .A(B[18]), .B(carry[18]), .Y(n5) );
  XOR2X1 U8 ( .A(B[18]), .B(carry[18]), .Y(SUM[18]) );
endmodule


module DPA_DW01_add_26 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [19:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U3 ( .A(A[19]), .B(carry[19]), .Y(SUM[19]) );
endmodule


module DPA_DW01_add_27 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [19:1] carry;

  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR2X1 U1 ( .A(A[17]), .B(n2), .Y(SUM[17]) );
  XOR2X1 U2 ( .A(A[16]), .B(n3), .Y(SUM[16]) );
  XOR2X1 U3 ( .A(A[15]), .B(n4), .Y(SUM[15]) );
  XOR2X1 U4 ( .A(A[14]), .B(n5), .Y(SUM[14]) );
  XOR2X1 U5 ( .A(A[13]), .B(n6), .Y(SUM[13]) );
  XOR2X1 U6 ( .A(A[12]), .B(n7), .Y(SUM[12]) );
  XOR2X1 U7 ( .A(A[11]), .B(n8), .Y(SUM[11]) );
  AND2X2 U8 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2X1 U9 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  AND2X2 U10 ( .A(A[16]), .B(n3), .Y(n2) );
  AND2X2 U11 ( .A(A[15]), .B(n4), .Y(n3) );
  AND2X2 U12 ( .A(A[14]), .B(n5), .Y(n4) );
  AND2X2 U13 ( .A(A[13]), .B(n6), .Y(n5) );
  AND2X2 U14 ( .A(A[12]), .B(n7), .Y(n6) );
  AND2X2 U15 ( .A(A[11]), .B(n8), .Y(n7) );
  AND2X2 U16 ( .A(A[10]), .B(carry[10]), .Y(n8) );
  CLKBUFX2 U17 ( .A(B[1]), .Y(SUM[1]) );
  CLKBUFX3 U18 ( .A(B[0]), .Y(SUM[0]) );
  AND2X2 U19 ( .A(A[17]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U20 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
endmodule


module DPA_DW01_add_28 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [19:1] carry;

  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U3 ( .A(A[17]), .B(n3), .Y(n2) );
  AND2X2 U4 ( .A(A[16]), .B(carry[16]), .Y(n3) );
  XNOR2X1 U5 ( .A(A[19]), .B(n4), .Y(SUM[19]) );
  NAND2X1 U6 ( .A(A[18]), .B(n2), .Y(n4) );
  XOR2X1 U7 ( .A(A[18]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U8 ( .A(A[17]), .B(n3), .Y(SUM[17]) );
  XOR2X1 U9 ( .A(A[16]), .B(carry[16]), .Y(SUM[16]) );
endmodule


module DPA_DW01_add_29 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [19:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X2 U2 ( .A(B[17]), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(B[16]), .B(carry[16]), .Y(n3) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X1 U5 ( .A(B[19]), .B(n4), .Y(SUM[19]) );
  NAND2X1 U6 ( .A(B[18]), .B(n2), .Y(n4) );
  XOR2X1 U7 ( .A(B[18]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U8 ( .A(B[17]), .B(n3), .Y(SUM[17]) );
  XOR2X1 U9 ( .A(B[16]), .B(carry[16]), .Y(SUM[16]) );
endmodule


module DPA_DW01_add_30 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [19:1] carry;

  CMPR32X2 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CMPR32X2 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(A[9]), .B(n12), .Y(SUM[9]) );
  XOR2X1 U2 ( .A(A[8]), .B(n13), .Y(SUM[8]) );
  CLKXOR2X2 U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X2 U5 ( .A(A[18]), .B(n3), .Y(n2) );
  XOR2X1 U6 ( .A(A[12]), .B(n9), .Y(SUM[12]) );
  XOR2X1 U7 ( .A(A[10]), .B(n11), .Y(SUM[10]) );
  XOR2X1 U8 ( .A(A[15]), .B(n6), .Y(SUM[15]) );
  XOR2X1 U9 ( .A(A[14]), .B(n7), .Y(SUM[14]) );
  XOR2X1 U10 ( .A(A[13]), .B(n8), .Y(SUM[13]) );
  XOR2X1 U11 ( .A(A[11]), .B(n10), .Y(SUM[11]) );
  XOR2X1 U12 ( .A(A[7]), .B(n14), .Y(SUM[7]) );
  XOR2X1 U13 ( .A(A[6]), .B(n15), .Y(SUM[6]) );
  XOR2X1 U14 ( .A(A[5]), .B(n16), .Y(SUM[5]) );
  AND2X2 U15 ( .A(A[17]), .B(n4), .Y(n3) );
  AND2X2 U16 ( .A(A[16]), .B(n5), .Y(n4) );
  AND2X2 U17 ( .A(A[15]), .B(n6), .Y(n5) );
  AND2X2 U18 ( .A(A[14]), .B(n7), .Y(n6) );
  AND2X2 U19 ( .A(A[13]), .B(n8), .Y(n7) );
  AND2X2 U20 ( .A(A[12]), .B(n9), .Y(n8) );
  AND2X2 U21 ( .A(A[11]), .B(n10), .Y(n9) );
  AND2X2 U22 ( .A(A[10]), .B(n11), .Y(n10) );
  AND2X2 U23 ( .A(A[9]), .B(n12), .Y(n11) );
  AND2X2 U24 ( .A(A[8]), .B(n13), .Y(n12) );
  AND2X2 U25 ( .A(A[7]), .B(n14), .Y(n13) );
  AND2X2 U26 ( .A(A[6]), .B(n15), .Y(n14) );
  AND2X2 U27 ( .A(A[5]), .B(n16), .Y(n15) );
  AND2X2 U28 ( .A(A[4]), .B(carry[4]), .Y(n16) );
  CLKXOR2X2 U29 ( .A(A[19]), .B(n2), .Y(SUM[19]) );
  CLKXOR2X2 U30 ( .A(A[18]), .B(n3), .Y(SUM[18]) );
  CLKXOR2X2 U31 ( .A(A[17]), .B(n4), .Y(SUM[17]) );
  CLKXOR2X2 U32 ( .A(A[16]), .B(n5), .Y(SUM[16]) );
  XOR2X1 U33 ( .A(A[4]), .B(carry[4]), .Y(SUM[4]) );
endmodule


module DPA_DW01_inc_6 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_80 ( A, B, CI, SUM, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [25:1] carry;

  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_79 ( A, B, CI, SUM, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [25:1] carry;

  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(SUM[25]), .S(
        SUM[24]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  OAI2BB1X1 U1 ( .A0N(A[1]), .A1N(B[1]), .B0(n1), .Y(carry[2]) );
  OAI211X1 U2 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n1) );
endmodule


module DPA_DW01_add_72 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   \carry[9] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n18;
  assign \carry[9]  = B[8];

  AND2XL U1 ( .A(B[9]), .B(\carry[9] ), .Y(n9) );
  AND2X2 U2 ( .A(B[17]), .B(n2), .Y(n1) );
  AND2X2 U3 ( .A(B[16]), .B(n3), .Y(n2) );
  AND2X2 U4 ( .A(B[15]), .B(n4), .Y(n3) );
  AND2X2 U5 ( .A(B[14]), .B(n5), .Y(n4) );
  AND2X2 U6 ( .A(B[13]), .B(n6), .Y(n5) );
  AND2X2 U7 ( .A(B[12]), .B(n7), .Y(n6) );
  AND2X2 U8 ( .A(B[11]), .B(n8), .Y(n7) );
  AND2X2 U9 ( .A(B[10]), .B(n9), .Y(n8) );
  NAND2XL U10 ( .A(B[18]), .B(n1), .Y(n18) );
  XOR2X1 U11 ( .A(B[18]), .B(n1), .Y(SUM[18]) );
  XOR2XL U12 ( .A(B[17]), .B(n2), .Y(SUM[17]) );
  XOR2XL U13 ( .A(B[16]), .B(n3), .Y(SUM[16]) );
  XOR2XL U14 ( .A(B[15]), .B(n4), .Y(SUM[15]) );
  XOR2XL U15 ( .A(B[14]), .B(n5), .Y(SUM[14]) );
  XOR2XL U16 ( .A(B[13]), .B(n6), .Y(SUM[13]) );
  XOR2XL U17 ( .A(B[12]), .B(n7), .Y(SUM[12]) );
  XOR2XL U18 ( .A(B[11]), .B(n8), .Y(SUM[11]) );
  XOR2XL U19 ( .A(B[10]), .B(n9), .Y(SUM[10]) );
  XOR2XL U20 ( .A(B[9]), .B(\carry[9] ), .Y(SUM[9]) );
  INVXL U21 ( .A(\carry[9] ), .Y(SUM[8]) );
  XNOR2X1 U22 ( .A(B[19]), .B(n18), .Y(SUM[19]) );
  CLKBUFX2 U23 ( .A(B[0]), .Y(SUM[0]) );
  CLKBUFX2 U24 ( .A(B[1]), .Y(SUM[1]) );
  CLKBUFX2 U25 ( .A(B[2]), .Y(SUM[2]) );
  CLKBUFX2 U26 ( .A(B[3]), .Y(SUM[3]) );
  CLKBUFX2 U27 ( .A(B[4]), .Y(SUM[4]) );
  CLKBUFX2 U28 ( .A(B[5]), .Y(SUM[5]) );
  CLKBUFX2 U29 ( .A(B[6]), .Y(SUM[6]) );
  CLKBUFX2 U30 ( .A(B[7]), .Y(SUM[7]) );
endmodule


module DPA_DW01_add_71 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n4;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  NAND2X1 U2 ( .A(A[18]), .B(carry[18]), .Y(n4) );
  XOR2X1 U3 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  XNOR2X1 U4 ( .A(A[19]), .B(n4), .Y(SUM[19]) );
  XOR2X1 U5 ( .A(A[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKBUFX3 U6 ( .A(A[0]), .Y(SUM[0]) );
  CLKBUFX3 U7 ( .A(A[1]), .Y(SUM[1]) );
endmodule


module DPA_DW01_add_70 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [19:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(A[19]), .B(carry[19]), .Y(SUM[19]) );
  XOR2XL U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_67 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n5;
  wire   [19:1] carry;

  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(n3) );
  AND2X2 U2 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2X1 U3 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  XNOR2X1 U4 ( .A(A[19]), .B(n5), .Y(SUM[19]) );
  NAND2X1 U5 ( .A(A[18]), .B(carry[18]), .Y(n5) );
  XOR2X1 U6 ( .A(A[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKINVX1 U7 ( .A(n3), .Y(SUM[0]) );
  CLKBUFX3 U8 ( .A(A[1]), .Y(SUM[1]) );
endmodule


module DPA_DW01_add_66 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;

  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  OR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[19]), .B(carry[19]), .Y(SUM[19]) );
  XNOR2XL U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_63 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  CLKBUFX3 U1 ( .A(B[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U3 ( .A(B[17]), .B(carry[17]), .Y(n2) );
  XOR2X1 U4 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  XNOR2X1 U5 ( .A(B[19]), .B(n4), .Y(SUM[19]) );
  NAND2X1 U6 ( .A(B[18]), .B(n2), .Y(n4) );
  XOR2X1 U7 ( .A(B[18]), .B(n2), .Y(SUM[18]) );
  XOR2XL U8 ( .A(B[17]), .B(carry[17]), .Y(SUM[17]) );
endmodule


module DPA_DW01_add_41 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n3;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  XNOR2X1 U3 ( .A(A[19]), .B(n3), .Y(SUM[19]) );
  NAND2X1 U4 ( .A(A[18]), .B(carry[18]), .Y(n3) );
  XOR2XL U5 ( .A(A[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKBUFX2 U6 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_74 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n3) );
  AND2X2 U2 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U3 ( .A(B[17]), .B(carry[17]), .Y(n2) );
  XOR2X1 U4 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  XNOR2X1 U5 ( .A(B[19]), .B(n5), .Y(SUM[19]) );
  NAND2X1 U6 ( .A(B[18]), .B(n2), .Y(n5) );
  XOR2X1 U7 ( .A(B[18]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U8 ( .A(B[17]), .B(carry[17]), .Y(SUM[17]) );
  CLKINVX1 U9 ( .A(n3), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_78 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [19:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X2 U2 ( .A(A[18]), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(A[17]), .B(n4), .Y(n3) );
  AND2X2 U4 ( .A(A[16]), .B(carry[16]), .Y(n4) );
  XOR2X1 U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XL U6 ( .A(A[19]), .B(n2), .Y(SUM[19]) );
  XOR2XL U7 ( .A(A[18]), .B(n3), .Y(SUM[18]) );
  XOR2XL U8 ( .A(A[17]), .B(n4), .Y(SUM[17]) );
  XOR2XL U9 ( .A(A[16]), .B(carry[16]), .Y(SUM[16]) );
endmodule


module DPA_DW01_add_77 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [19:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  XOR3X1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .Y(SUM[19]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_75 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n3;
  wire   [19:1] carry;
  assign carry[2] = B[1];

  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n1) );
  CLKINVX1 U2 ( .A(carry[2]), .Y(SUM[1]) );
  CLKINVX1 U3 ( .A(n1), .Y(SUM[0]) );
  XNOR2X1 U4 ( .A(B[19]), .B(n3), .Y(SUM[19]) );
  NAND2X1 U5 ( .A(B[18]), .B(carry[18]), .Y(n3) );
  XOR2X1 U6 ( .A(B[18]), .B(carry[18]), .Y(SUM[18]) );
endmodule


module DPA_DW01_add_44 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16;
  wire   [19:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U2 ( .A(B[17]), .B(n3), .Y(n2) );
  NAND2XL U3 ( .A(B[18]), .B(n2), .Y(n16) );
  XOR2X1 U4 ( .A(B[18]), .B(n2), .Y(SUM[18]) );
  AND2X2 U5 ( .A(B[16]), .B(n4), .Y(n3) );
  AND2X2 U6 ( .A(B[15]), .B(n5), .Y(n4) );
  AND2X2 U7 ( .A(B[14]), .B(n6), .Y(n5) );
  AND2X2 U8 ( .A(B[13]), .B(n7), .Y(n6) );
  AND2X2 U9 ( .A(B[12]), .B(n8), .Y(n7) );
  AND2X2 U10 ( .A(B[11]), .B(n9), .Y(n8) );
  AND2X2 U11 ( .A(B[10]), .B(n10), .Y(n9) );
  AND2X2 U12 ( .A(B[9]), .B(n11), .Y(n10) );
  AND2X2 U13 ( .A(B[8]), .B(n12), .Y(n11) );
  AND2X2 U14 ( .A(B[7]), .B(n13), .Y(n12) );
  AND2X2 U15 ( .A(B[6]), .B(n14), .Y(n13) );
  AND2X2 U16 ( .A(B[5]), .B(carry[5]), .Y(n14) );
  XNOR2X1 U17 ( .A(B[19]), .B(n16), .Y(SUM[19]) );
  XOR2XL U18 ( .A(B[17]), .B(n3), .Y(SUM[17]) );
  XOR2XL U19 ( .A(B[16]), .B(n4), .Y(SUM[16]) );
  XOR2XL U20 ( .A(B[15]), .B(n5), .Y(SUM[15]) );
  XOR2XL U21 ( .A(B[14]), .B(n6), .Y(SUM[14]) );
  XOR2XL U22 ( .A(B[13]), .B(n7), .Y(SUM[13]) );
  XOR2XL U23 ( .A(B[12]), .B(n8), .Y(SUM[12]) );
  XOR2XL U24 ( .A(B[11]), .B(n9), .Y(SUM[11]) );
  XOR2XL U25 ( .A(B[10]), .B(n10), .Y(SUM[10]) );
  XOR2XL U26 ( .A(B[9]), .B(n11), .Y(SUM[9]) );
  XOR2XL U27 ( .A(B[8]), .B(n12), .Y(SUM[8]) );
  XOR2XL U28 ( .A(B[7]), .B(n13), .Y(SUM[7]) );
  XOR2XL U29 ( .A(B[6]), .B(n14), .Y(SUM[6]) );
  XOR2XL U30 ( .A(B[5]), .B(carry[5]), .Y(SUM[5]) );
  XOR2XL U31 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
  CLKBUFX2 U32 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_43 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n4;
  wire   [19:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  NAND2X1 U2 ( .A(B[18]), .B(carry[18]), .Y(n4) );
  XNOR2X1 U3 ( .A(B[19]), .B(n4), .Y(SUM[19]) );
  XOR2X1 U4 ( .A(B[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKBUFX2 U5 ( .A(B[1]), .Y(SUM[1]) );
  CLKBUFX3 U6 ( .A(B[0]), .Y(SUM[0]) );
  XOR2XL U7 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
endmodule


module DPA_DW01_add_33 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_32 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_31 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [10:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(SUM[9]), .S(SUM[8]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  OAI2BB1X1 U1 ( .A0N(A[1]), .A1N(B[1]), .B0(n1), .Y(carry[2]) );
  OAI211X1 U2 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n1) );
endmodule


module DPA_DW01_add_46 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [19:1] carry;
  assign carry[1] = B[0];

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[17]), .B(n2), .Y(n1) );
  NAND2XL U2 ( .A(B[18]), .B(n1), .Y(n14) );
  XOR2X1 U3 ( .A(B[18]), .B(n1), .Y(SUM[18]) );
  AND2X2 U4 ( .A(B[16]), .B(n3), .Y(n2) );
  AND2X2 U5 ( .A(B[15]), .B(n4), .Y(n3) );
  AND2X2 U6 ( .A(B[14]), .B(n5), .Y(n4) );
  AND2X2 U7 ( .A(B[13]), .B(n6), .Y(n5) );
  AND2X2 U8 ( .A(B[12]), .B(n7), .Y(n6) );
  AND2X2 U9 ( .A(B[11]), .B(n8), .Y(n7) );
  AND2X2 U10 ( .A(B[10]), .B(n9), .Y(n8) );
  AND2X2 U11 ( .A(B[9]), .B(n10), .Y(n9) );
  AND2X2 U12 ( .A(B[8]), .B(n11), .Y(n10) );
  AND2X2 U13 ( .A(B[7]), .B(n12), .Y(n11) );
  AND2X2 U14 ( .A(B[6]), .B(n13), .Y(n12) );
  AND2X2 U15 ( .A(B[5]), .B(carry[5]), .Y(n13) );
  XNOR2X1 U16 ( .A(B[19]), .B(n14), .Y(SUM[19]) );
  XOR2XL U17 ( .A(B[17]), .B(n2), .Y(SUM[17]) );
  XOR2XL U18 ( .A(B[16]), .B(n3), .Y(SUM[16]) );
  XOR2XL U19 ( .A(B[15]), .B(n4), .Y(SUM[15]) );
  XOR2XL U20 ( .A(B[14]), .B(n5), .Y(SUM[14]) );
  XOR2XL U21 ( .A(B[13]), .B(n6), .Y(SUM[13]) );
  XOR2XL U22 ( .A(B[12]), .B(n7), .Y(SUM[12]) );
  XOR2XL U23 ( .A(B[11]), .B(n8), .Y(SUM[11]) );
  XOR2XL U24 ( .A(B[10]), .B(n9), .Y(SUM[10]) );
  XOR2XL U25 ( .A(B[9]), .B(n10), .Y(SUM[9]) );
  XOR2XL U26 ( .A(B[8]), .B(n11), .Y(SUM[8]) );
  XOR2XL U27 ( .A(B[7]), .B(n12), .Y(SUM[7]) );
  XOR2XL U28 ( .A(B[6]), .B(n13), .Y(SUM[6]) );
  XOR2XL U29 ( .A(B[5]), .B(carry[5]), .Y(SUM[5]) );
  CLKINVX1 U30 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_45 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n4;
  wire   [19:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  NAND2X1 U2 ( .A(B[18]), .B(carry[18]), .Y(n4) );
  XNOR2X1 U3 ( .A(B[19]), .B(n4), .Y(SUM[19]) );
  XOR2X1 U4 ( .A(B[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKBUFX3 U5 ( .A(B[0]), .Y(SUM[0]) );
  XOR2XL U6 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U7 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module DPA_DW01_add_48 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [19:1] carry;
  assign carry[1] = B[0];

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[17]), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(B[16]), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(B[15]), .B(n4), .Y(n3) );
  AND2X2 U4 ( .A(B[14]), .B(n5), .Y(n4) );
  AND2X2 U5 ( .A(B[13]), .B(n6), .Y(n5) );
  AND2X2 U6 ( .A(B[12]), .B(n7), .Y(n6) );
  AND2X2 U7 ( .A(B[11]), .B(n8), .Y(n7) );
  AND2X2 U8 ( .A(B[10]), .B(n9), .Y(n8) );
  AND2X2 U9 ( .A(B[9]), .B(n10), .Y(n9) );
  AND2X2 U10 ( .A(B[8]), .B(n11), .Y(n10) );
  AND2X2 U11 ( .A(B[7]), .B(n12), .Y(n11) );
  AND2X2 U12 ( .A(B[6]), .B(n13), .Y(n12) );
  AND2X2 U13 ( .A(B[5]), .B(carry[5]), .Y(n13) );
  AND2X2 U14 ( .A(B[18]), .B(n1), .Y(n14) );
  XOR2X1 U15 ( .A(B[18]), .B(n1), .Y(SUM[18]) );
  XOR2XL U16 ( .A(B[17]), .B(n2), .Y(SUM[17]) );
  XOR2XL U17 ( .A(B[16]), .B(n3), .Y(SUM[16]) );
  XOR2XL U18 ( .A(B[15]), .B(n4), .Y(SUM[15]) );
  XOR2XL U19 ( .A(B[14]), .B(n5), .Y(SUM[14]) );
  XOR2XL U20 ( .A(B[13]), .B(n6), .Y(SUM[13]) );
  XOR2XL U21 ( .A(B[12]), .B(n7), .Y(SUM[12]) );
  XOR2XL U22 ( .A(B[11]), .B(n8), .Y(SUM[11]) );
  XOR2XL U23 ( .A(B[10]), .B(n9), .Y(SUM[10]) );
  XOR2XL U24 ( .A(B[9]), .B(n10), .Y(SUM[9]) );
  XOR2XL U25 ( .A(B[8]), .B(n11), .Y(SUM[8]) );
  XOR2XL U26 ( .A(B[7]), .B(n12), .Y(SUM[7]) );
  XOR2XL U27 ( .A(B[6]), .B(n13), .Y(SUM[6]) );
  XOR2XL U28 ( .A(B[5]), .B(carry[5]), .Y(SUM[5]) );
  XOR2XL U29 ( .A(B[19]), .B(n14), .Y(SUM[19]) );
  CLKINVX1 U30 ( .A(carry[1]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_47 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  AND2X2 U2 ( .A(B[18]), .B(carry[18]), .Y(n2) );
  XOR2XL U3 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  XOR2X1 U4 ( .A(B[19]), .B(n2), .Y(SUM[19]) );
  XOR2X1 U5 ( .A(B[18]), .B(carry[18]), .Y(SUM[18]) );
  CLKBUFX3 U6 ( .A(B[1]), .Y(SUM[1]) );
  CLKBUFX3 U7 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_51 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [19:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X2 U2 ( .A(B[18]), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(B[17]), .B(n4), .Y(n3) );
  AND2X2 U4 ( .A(B[16]), .B(n5), .Y(n4) );
  AND2X2 U5 ( .A(B[15]), .B(n6), .Y(n5) );
  AND2X2 U6 ( .A(B[14]), .B(n7), .Y(n6) );
  AND2X2 U7 ( .A(B[13]), .B(n8), .Y(n7) );
  AND2X2 U8 ( .A(B[12]), .B(n9), .Y(n8) );
  AND2X2 U9 ( .A(B[11]), .B(n10), .Y(n9) );
  AND2X2 U10 ( .A(B[10]), .B(n11), .Y(n10) );
  AND2X2 U11 ( .A(B[9]), .B(n12), .Y(n11) );
  AND2X2 U12 ( .A(B[8]), .B(carry[8]), .Y(n12) );
  XOR2XL U13 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XL U14 ( .A(B[19]), .B(n2), .Y(SUM[19]) );
  XOR2X1 U15 ( .A(B[18]), .B(n3), .Y(SUM[18]) );
  XOR2X1 U16 ( .A(B[17]), .B(n4), .Y(SUM[17]) );
  XOR2XL U17 ( .A(B[16]), .B(n5), .Y(SUM[16]) );
  XOR2XL U18 ( .A(B[15]), .B(n6), .Y(SUM[15]) );
  XOR2XL U19 ( .A(B[14]), .B(n7), .Y(SUM[14]) );
  XOR2XL U20 ( .A(B[13]), .B(n8), .Y(SUM[13]) );
  XOR2XL U21 ( .A(B[12]), .B(n9), .Y(SUM[12]) );
  XOR2XL U22 ( .A(B[11]), .B(n10), .Y(SUM[11]) );
  XOR2XL U23 ( .A(B[10]), .B(n11), .Y(SUM[10]) );
  XOR2XL U24 ( .A(B[9]), .B(n12), .Y(SUM[9]) );
  XOR2XL U25 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module DPA_DW01_add_50 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [19:1] carry;

  AND2X2 U1 ( .A(B[18]), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(B[17]), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(B[16]), .B(carry[16]), .Y(n3) );
  OR2X1 U4 ( .A(B[15]), .B(carry[15]), .Y(carry[16]) );
  OR2X1 U5 ( .A(B[14]), .B(carry[14]), .Y(carry[15]) );
  OR2X1 U6 ( .A(B[13]), .B(n4), .Y(carry[14]) );
  AND2X2 U7 ( .A(B[12]), .B(carry[12]), .Y(n4) );
  OR2X1 U8 ( .A(B[11]), .B(n5), .Y(carry[12]) );
  AND2X2 U9 ( .A(B[10]), .B(n6), .Y(n5) );
  AND2X2 U10 ( .A(B[9]), .B(n7), .Y(n6) );
  AND2X2 U11 ( .A(B[8]), .B(A[8]), .Y(n7) );
  XOR2X1 U12 ( .A(B[19]), .B(n1), .Y(SUM[19]) );
  XOR2X1 U13 ( .A(B[18]), .B(n2), .Y(SUM[18]) );
  XOR2X1 U14 ( .A(B[17]), .B(n3), .Y(SUM[17]) );
  XOR2X1 U15 ( .A(B[16]), .B(carry[16]), .Y(SUM[16]) );
  XNOR2X1 U16 ( .A(B[15]), .B(carry[15]), .Y(SUM[15]) );
  XNOR2X1 U17 ( .A(B[14]), .B(carry[14]), .Y(SUM[14]) );
  XNOR2X1 U18 ( .A(B[13]), .B(n4), .Y(SUM[13]) );
  XOR2X1 U19 ( .A(B[12]), .B(carry[12]), .Y(SUM[12]) );
  XNOR2X1 U20 ( .A(B[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U21 ( .A(B[10]), .B(n6), .Y(SUM[10]) );
  XOR2X1 U22 ( .A(B[9]), .B(n7), .Y(SUM[9]) );
  XOR2X1 U23 ( .A(B[8]), .B(A[8]), .Y(SUM[8]) );
  CLKBUFX3 U24 ( .A(A[7]), .Y(SUM[7]) );
  CLKBUFX3 U25 ( .A(A[6]), .Y(SUM[6]) );
  CLKBUFX3 U26 ( .A(A[5]), .Y(SUM[5]) );
  CLKBUFX3 U27 ( .A(A[4]), .Y(SUM[4]) );
  CLKBUFX3 U28 ( .A(A[3]), .Y(SUM[3]) );
  CLKBUFX3 U29 ( .A(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U30 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U31 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DPA_DW01_add_49 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [19:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  XOR3X1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .Y(SUM[19]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module DPA ( clk, reset, IM_A, IM_Q, IM_D, IM_WEN, CR_A, CR_Q );
  output [19:0] IM_A;
  input [23:0] IM_Q;
  output [23:0] IM_D;
  output [8:0] CR_A;
  input [12:0] CR_Q;
  input clk, reset;
  output IM_WEN;
  wire   n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, \IM_D_t[0][23] ,
         \IM_D_t[0][22] , \IM_D_t[0][21] , \IM_D_t[0][20] , \IM_D_t[0][19] ,
         \IM_D_t[0][18] , \IM_D_t[0][17] , \IM_D_t[0][16] , \IM_D_t[0][15] ,
         \IM_D_t[0][14] , \IM_D_t[0][13] , \IM_D_t[0][12] , \IM_D_t[0][11] ,
         \IM_D_t[0][10] , \IM_D_t[0][9] , \IM_D_t[0][8] , \IM_D_t[0][7] ,
         \IM_D_t[0][6] , \IM_D_t[0][5] , \IM_D_t[0][4] , \IM_D_t[0][3] ,
         \IM_D_t[0][2] , \IM_D_t[0][1] , \IM_D_t[0][0] , \IM_D_t[1][23] ,
         \IM_D_t[1][22] , \IM_D_t[1][21] , \IM_D_t[1][20] , \IM_D_t[1][19] ,
         \IM_D_t[1][18] , \IM_D_t[1][17] , \IM_D_t[1][16] , \IM_D_t[1][15] ,
         \IM_D_t[1][14] , \IM_D_t[1][13] , \IM_D_t[1][12] , \IM_D_t[1][11] ,
         \IM_D_t[1][10] , \IM_D_t[1][9] , \IM_D_t[1][8] , \IM_D_t[1][7] ,
         \IM_D_t[1][6] , \IM_D_t[1][5] , \IM_D_t[1][4] , \IM_D_t[1][3] ,
         \IM_D_t[1][2] , \IM_D_t[1][1] , \IM_D_t[1][0] , \IM_D_t[2][23] ,
         \IM_D_t[2][22] , \IM_D_t[2][21] , \IM_D_t[2][20] , \IM_D_t[2][19] ,
         \IM_D_t[2][18] , \IM_D_t[2][17] , \IM_D_t[2][16] , \IM_D_t[2][15] ,
         \IM_D_t[2][14] , \IM_D_t[2][13] , \IM_D_t[2][12] , \IM_D_t[2][11] ,
         \IM_D_t[2][10] , \IM_D_t[2][9] , \IM_D_t[2][8] , \IM_D_t[2][7] ,
         \IM_D_t[2][6] , \IM_D_t[2][5] , \IM_D_t[2][4] , \IM_D_t[2][3] ,
         \IM_D_t[2][2] , \IM_D_t[2][1] , \IM_D_t[2][0] , \IM_D_t[3][23] ,
         \IM_D_t[3][22] , \IM_D_t[3][21] , \IM_D_t[3][20] , \IM_D_t[3][19] ,
         \IM_D_t[3][18] , \IM_D_t[3][17] , \IM_D_t[3][16] , \IM_D_t[3][15] ,
         \IM_D_t[3][14] , \IM_D_t[3][13] , \IM_D_t[3][12] , \IM_D_t[3][11] ,
         \IM_D_t[3][10] , \IM_D_t[3][9] , \IM_D_t[3][8] , \IM_D_t[3][7] ,
         \IM_D_t[3][6] , \IM_D_t[3][5] , \IM_D_t[3][4] , \IM_D_t[3][3] ,
         \IM_D_t[3][2] , \IM_D_t[3][1] , \IM_D_t[3][0] , N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N444,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477,
         N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N501, N502, N503, N504, N505, N506, N508, N509, N510, N511,
         N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522,
         N523, N524, N525, N526, N527, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564,
         N565, N566, N567, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698,
         N699, N700, N701, N702, N703, N704, N705, N706, N707, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, N727, N728, N807, N808, N809, N810,
         N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821,
         N822, N823, N824, N825, N826, N867, N868, N869, N870, N871, N872,
         N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883,
         N884, N885, N886, N944, N945, N946, N947, N948, N949, N950, N951,
         N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962,
         N963, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032,
         N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042,
         N1043, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287,
         N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297,
         N1298, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364,
         N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374,
         N1375, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449,
         N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459,
         N1460, N2136, N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189,
         N2190, N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199,
         N2200, N2201, N2202, N2203, N2204, N2205, N2318, N2319, N2320, N2321,
         N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331,
         N2332, N2333, N2334, N2335, N2336, N2337, N2413, N2414, N2415, N2416,
         N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2488, N2489, N2490,
         N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500,
         N2501, N2502, N2503, N2785, N2786, N2787, N2788, N2789, N2790, N2791,
         N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799, N2800, N2801,
         N2802, N2803, N2804, N2850, N2851, N2852, N2853, N2854, N2855, N2856,
         N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866,
         N2867, N2868, N2869, N2944, N2945, N2946, N2947, N2948, N2949, N2950,
         N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2984,
         N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994,
         N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004,
         N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3213, N3214,
         N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224,
         N3225, N3226, N3227, N3228, N3617, N3618, N3619, N3620, N3621, N3622,
         N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632,
         N3633, N3634, N3635, N3636, N3662, N3663, N3664, N3665, N3666, N3667,
         N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677,
         N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3688,
         N3689, N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698,
         N3699, N3700, N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708,
         N3709, N3710, N3711, N3732, N3733, N3734, N3735, N3736, N3737, N3738,
         N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748,
         N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758,
         N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768,
         N3769, N3770, N3771, N3841, N4086, N4087, N4088, N4089, N4090, N4091,
         N4092, N4093, N4094, N4095, N4096, N4097, N4098, N4099, N4100, N4101,
         N4102, N4103, N4104, N4105, N4106, N4107, N4108, N4109, N4110, N4111,
         N4112, N4113, N4114, N4115, N4116, N4117, N4118, N4119, N4120, N4121,
         N4122, N4123, N4124, N4125, N4176, N4177, N4178, N4179, N4180, N4181,
         N4182, N4183, N4184, N4185, N4186, N4187, N4188, N4189, N4190, N4191,
         N4192, N4193, N4194, N4195, N4271, N4272, N4273, N4274, N4275, N4276,
         N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284, N4285, N4286,
         N4287, N4288, N4289, N4290, N4291, N4292, N4293, N4294, N4364, N4365,
         N4366, N4367, N4368, N4369, N4370, N4371, N4372, N4373, N4374, N4375,
         N4376, N4377, N4378, N4379, N4380, N4381, N4382, N4383, N4409, N4410,
         N4411, N4412, N4413, N4414, N4415, N4416, N4417, N4418, N4419, N4420,
         N4421, N4422, N4423, N4424, N4425, N4426, N4427, N4428, N4454, N4455,
         N4456, N4457, N4458, N4459, N4460, N4461, N4462, N4463, N4464, N4465,
         N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473, N4615, N4616,
         N4617, N4618, N4619, N4620, N4621, N4622, N4623, N4624, N4625, N4626,
         N4627, N4628, N4629, N4630, N4631, N4632, N4633, N4634, N4635, N4636,
         N4637, N4638, N4639, N4640, N4641, N4642, N4643, N4644, N4645, N4646,
         N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985,
         N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994, N4995,
         N5021, N5022, N5023, N5024, N5025, N5026, N5027, N5028, N5029, N5030,
         N5031, N5032, N5033, N5034, N5035, N5036, N5037, N5038, N5039, N5040,
         N5147, N5148, N5149, N5150, N5151, N5152, N5153, N5154, N5155, N5156,
         N5157, N5158, N5159, N5160, N5161, N5162, N5163, N5164, N5165, N5166,
         N5167, N5852, N5853, N5854, N5855, N5856, N5862, N5863, N5864, N5865,
         N5892, N5893, N5894, N5895, N5896, N5897, N5919, N5920, N5921, N5922,
         N5923, N5924, N5945, N5946, N5947, N5948, N5949, N5950, N5965, N5966,
         N5967, N5968, N6005, N6006, N6007, N6008, N6009, N6017, N6018, N6019,
         N6024, N6025, N6026, N6027, N6028, N6061, N6062, N6063, N6064, N6065,
         N6066, N6088, N6089, N6090, N6091, N6092, N6093, N6115, N6116, N6117,
         N6118, N6119, N6120, N6142, N6143, N6144, N6145, N6146, N6147, N6169,
         N6170, N6171, N6172, N6173, N6174, N6195, N6196, N6197, N6198, N6199,
         N6200, N6302, N6303, N6304, N6305, N6306, N6307, N6329, N6330, N6331,
         N6332, N6333, N6334, N6356, N6357, N6358, N6359, N6360, N6361, N6383,
         N6384, N6385, N6386, N6387, N6388, N6410, N6411, N6412, N6413, N6414,
         N6415, N6436, N6437, N6438, N6439, N6440, N6441, N6550, N6551, N6552,
         N6553, N6554, N6555, N6556, N6557, N6558, N6559, N6560, N6561, N6562,
         N6563, N6564, N6565, N6566, N6567, N6568, N6569, N6745, N6746, N6747,
         N6748, N6749, N6750, N6751, N6752, N6753, N6754, N6755, N6756, N6757,
         N6758, N6759, N6760, N6761, N6762, N6763, N6764, N6769, N6770, N6771,
         N6772, N6773, N6774, N6775, N6783, N6784, N6785, N6786, N6787, N6788,
         N6789, N6804, N6805, N6806, N6807, N6808, N6809, N6810, N7625, N7626,
         N7627, N7628, N7629, N7630, N7631, N7632, N7633, N7634, N7635, N7636,
         N7637, N7638, N7639, N7640, N7641, N7642, N7643, N7644, N7645, N7646,
         N7647, N7648, N7649, N7650, N7651, N7652, N7653, N7654, N7655, N7656,
         N7657, N7658, N7659, N7660, N7661, N7662, N7663, N7664, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n137, n138, n139, n140, n141, n142, n143, n144,
         \gt_332/n15 , \gt_332/n9 , n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1927, n2016, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2098, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, N6165, N6164, N6163, N6162, N6161, N6160, N6154,
         N6153, N6151, N6150, N6406, N6405, N6404, N6403, N6402, N6401, N6395,
         N6394, N6392, N6391, N6191, N6190, N6189, N6188, N6187, N6180, N6179,
         N6178, N6177, N6138, N6137, N6136, N6135, N6134, N6127, N6126, N6125,
         N6124, N6432, N6431, N6430, N6429, N6428, N6421, N6420, N6419, N6418,
         N6379, N6378, N6377, N6376, N6375, N6368, N6367, N6366, N6365, N7684,
         N7683, N7682, N7681, N7680, N7679, N7678, N7677, N7676, N7675, N7674,
         N7673, N7672, N7671, N7670, N7669, N7668, N7667, N7666, N7622, N7621,
         N7620, N7619, N7618, N7617, N7616, N7615, N7614, N7613, N7612, N7611,
         N7610, N7609, N7608, N7607, N7606, N7605, N7604, N688, N687, N686,
         N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675,
         N674, N673, N672, N671, N670, N668, N667, N666, N2849, N2848, N2847,
         N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837,
         N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827,
         N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817,
         N2816, N2815, N2814, N2813, N2812, N2811, N1400, N1399, N1398, N1397,
         N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387,
         N1386, N1385, N1384, N1383, N1382, N4360, N4359, N4358, N4357, N4356,
         N4355, N4354, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345,
         N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334,
         N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4323,
         N4322, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696,
         N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686,
         N4433, N4432, N4431, N4429, N6111, N6110, N6109, N6108, N6107, N6100,
         N6099, N6098, N6352, N6351, N6350, N6349, N6348, N6341, N6340, N6339,
         N5915, N5914, N5913, N5912, N5911, N5910, N5904, N5903, N5902, N5901,
         N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269,
         N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259,
         N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1239, N804,
         N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793,
         N791, N790, N789, N6084, N6083, N6082, N6081, N6080, N6073, N6072,
         N6071, N6070, N6325, N6324, N6323, N6322, N6321, N6314, N6313, N6312,
         N6311, N5941, N5940, N5939, N5938, N5937, N5930, N5929, N5928, N5926,
         N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346,
         N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336,
         N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N623,
         N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612,
         N611, N610, N609, N608, N607, N606, N605, N604, N2764, N2763, N2762,
         N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752,
         N2751, N2750, N2749, N2748, N2747, N2746, N2745, N5888, N5887, N5886,
         N5885, N5884, N6549, N6548, N6547, N6546, N6545, N6544, N6543, N6542,
         N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534, N6533, N6532,
         N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524, N6523, N6522,
         N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514, N6513, N6512,
         N6511, N6510, N6509, N6508, N6507, N6506, N6505, N6504, N6490, N6489,
         N6488, N6487, N6486, N6484, N6483, N6482, N6057, N6056, N6055, N6054,
         N6053, N6298, N6297, N6296, N6295, N6294, \add_772/carry[6] ,
         \add_772/carry[7] , \add_772/carry[8] , \r1795/carry[5] ,
         \r1795/carry[6] , \r1795/carry[7] , \r1794/carry[7] ,
         \r1793/carry[7] , \r1778/carry[6] , \r1777/carry[5] ,
         \add_817/carry[8] , \add_817/carry[7] , \add_817/carry[6] ,
         \add_817/carry[5] , \mult_817/n5 , \mult_817/n4 , \mult_817/n3 ,
         \mult_817/n2 , \add_819/carry[8] , \add_819/carry[7] ,
         \add_819/carry[6] , \add_819/carry[5] , \mult_819/n5 , \mult_819/n4 ,
         \mult_819/n3 , \mult_819/n2 , \sub_819/carry[3] , \sub_819/carry[5] ,
         \add_821/carry[8] , \add_821/carry[7] , \add_821/carry[6] ,
         \add_821/carry[5] , \mult_821/n5 , \mult_821/n4 , \mult_821/n3 ,
         \mult_821/n2 , \sub_821/carry[4] , \add_823/carry[8] ,
         \add_823/carry[7] , \add_823/carry[6] , \add_823/carry[5] ,
         \mult_823/n5 , \mult_823/n4 , \mult_823/n3 , \mult_823/n2 ,
         \add_827/carry[8] , \add_827/carry[7] , \add_827/carry[6] ,
         \add_827/carry[5] , \mult_827/n5 , \mult_827/n4 , \mult_827/n3 ,
         \mult_827/n2 , \sub_827/carry[3] , \sub_827/carry[4] ,
         \add_825/carry[8] , \add_825/carry[7] , \add_825/carry[6] ,
         \add_825/carry[5] , \mult_825/n5 , \mult_825/n4 , \mult_825/n3 ,
         \mult_825/n2 , \sub_825/carry[5] ,
         \add_0_root_add_0_root_add_601_3/carry[19] ,
         \add_0_root_add_0_root_add_601_3/carry[18] ,
         \add_0_root_add_0_root_add_601_3/carry[17] ,
         \add_0_root_add_0_root_add_601_3/carry[16] ,
         \add_0_root_add_0_root_add_601_3/carry[15] ,
         \add_0_root_add_0_root_add_601_3/carry[14] ,
         \add_0_root_add_0_root_add_601_3/carry[13] ,
         \add_0_root_add_0_root_add_601_3/carry[12] ,
         \add_0_root_add_0_root_add_601_3/carry[11] ,
         \add_0_root_add_0_root_add_601_3/carry[10] ,
         \add_0_root_add_0_root_add_601_3/carry[9] ,
         \add_0_root_add_0_root_add_601_3/carry[8] ,
         \add_0_root_add_0_root_add_601_3/carry[7] ,
         \add_0_root_add_0_root_add_601_3/carry[6] ,
         \add_0_root_add_0_root_add_601_3/carry[5] ,
         \add_0_root_add_0_root_add_601_3/carry[4] ,
         \add_0_root_add_0_root_add_601_3/carry[3] , \sub_601/carry[4] ,
         \mult_869/n11 , \mult_869/n10 , \mult_869/n9 , \mult_869/n8 ,
         \mult_869/n7 , \mult_869/n6 , \mult_869/n5 , \mult_869/n4 ,
         \mult_869/n3 , \mult_869/n2 ,
         \add_3_root_add_0_root_add_869_4/carry[5] , \add_765/carry[8] ,
         \add_765/carry[7] , \add_765/carry[6] , \add_765/carry[5] ,
         \mult_765/n5 , \mult_765/n4 , \mult_765/n3 , \mult_765/n2 ,
         \add_769/carry[8] , \add_769/carry[7] , \add_769/carry[6] ,
         \add_769/carry[5] , \mult_769/n5 , \mult_769/n4 , \mult_769/n3 ,
         \mult_769/n2 , \sub_769/carry[4] , \add_767/carry[8] ,
         \add_767/carry[7] , \add_767/carry[6] , \add_767/carry[5] ,
         \mult_767/n5 , \mult_767/n4 , \mult_767/n3 , \mult_767/n2 ,
         \sub_767/carry[3] , \sub_767/carry[5] , \add_789/carry[8] ,
         \add_789/carry[7] , \add_789/carry[6] , \add_789/carry[5] ,
         \mult_789/n5 , \mult_789/n4 , \mult_789/n3 , \mult_789/n2 ,
         \add_791/carry[8] , \add_791/carry[7] , \add_791/carry[6] ,
         \add_791/carry[5] , \mult_791/n5 , \mult_791/n4 , \mult_791/n3 ,
         \mult_791/n2 , \sub_791/carry[3] , \sub_791/carry[5] ,
         \add_793/carry[8] , \add_793/carry[7] , \add_793/carry[6] ,
         \add_793/carry[5] , \mult_793/n5 , \mult_793/n4 , \mult_793/n3 ,
         \mult_793/n2 , \sub_793/carry[4] , \add_795/carry[8] ,
         \add_795/carry[7] , \add_795/carry[6] , \add_795/carry[5] ,
         \mult_795/n5 , \mult_795/n4 , \mult_795/n3 , \mult_795/n2 ,
         \add_799/carry[8] , \add_799/carry[7] , \add_799/carry[6] ,
         \add_799/carry[5] , \mult_799/n5 , \mult_799/n4 , \mult_799/n3 ,
         \mult_799/n2 , \sub_799/carry[3] , \sub_799/carry[4] ,
         \add_797/carry[8] , \add_797/carry[7] , \add_797/carry[6] ,
         \add_797/carry[5] , \mult_797/n5 , \mult_797/n4 , \mult_797/n3 ,
         \mult_797/n2 , \sub_797/carry[5] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[19] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[18] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[17] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[16] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[15] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[14] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[13] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[12] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[11] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[10] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[9] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[8] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[7] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[6] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[5] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[4] ,
         \add_0_root_add_0_root_add_579_4_cf/carry[3] ,
         \add_0_root_add_1_root_add_282_4/carry[19] ,
         \add_0_root_add_1_root_add_282_4/carry[18] ,
         \add_0_root_add_1_root_add_282_4/carry[17] ,
         \add_0_root_add_1_root_add_282_4/carry[16] ,
         \add_0_root_add_1_root_add_282_4/carry[15] ,
         \add_0_root_add_1_root_add_282_4/carry[14] ,
         \add_0_root_add_1_root_add_282_4/carry[13] ,
         \add_0_root_add_1_root_add_282_4/carry[12] ,
         \add_0_root_add_1_root_add_282_4/carry[11] ,
         \add_0_root_add_1_root_add_282_4/carry[10] ,
         \add_0_root_add_1_root_add_282_4/carry[9] ,
         \add_0_root_add_1_root_add_282_4/carry[8] ,
         \add_0_root_add_1_root_add_282_4/carry[7] ,
         \add_0_root_add_1_root_add_282_4/carry[6] ,
         \add_0_root_add_1_root_add_282_4/carry[5] ,
         \add_0_root_add_1_root_add_282_4/carry[4] ,
         \add_0_root_add_1_root_add_282_4/carry[3] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[19] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[18] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[17] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[16] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[15] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[14] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[13] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[12] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[11] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[10] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[9] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[8] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[7] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[6] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[5] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[4] ,
         \add_0_root_add_0_root_add_661_4_cf/carry[3] ,
         \add_0_root_add_0_root_add_209_3/carry[19] ,
         \add_0_root_add_0_root_add_209_3/carry[18] ,
         \add_0_root_add_0_root_add_209_3/carry[17] ,
         \add_0_root_add_0_root_add_209_3/carry[16] ,
         \add_0_root_add_0_root_add_209_3/carry[15] ,
         \add_0_root_add_0_root_add_209_3/carry[14] ,
         \add_0_root_add_0_root_add_209_3/carry[13] ,
         \add_0_root_add_0_root_add_209_3/carry[12] ,
         \add_0_root_add_0_root_add_209_3/carry[11] ,
         \add_0_root_add_0_root_add_209_3/carry[10] ,
         \add_0_root_add_0_root_add_209_3/carry[9] ,
         \add_0_root_add_0_root_add_209_3/carry[8] ,
         \add_0_root_add_0_root_add_209_3/carry[7] ,
         \add_0_root_add_0_root_add_209_3/carry[6] ,
         \add_0_root_add_0_root_add_209_3/carry[5] ,
         \add_0_root_add_0_root_add_209_3/carry[4] ,
         \add_0_root_add_0_root_add_209_3/carry[3] ,
         \add_0_root_add_0_root_add_446_3/carry[19] ,
         \add_0_root_add_0_root_add_446_3/carry[18] ,
         \add_0_root_add_0_root_add_446_3/carry[17] ,
         \add_0_root_add_0_root_add_446_3/carry[16] ,
         \add_0_root_add_0_root_add_446_3/carry[15] ,
         \add_0_root_add_0_root_add_446_3/carry[14] ,
         \add_0_root_add_0_root_add_446_3/carry[13] ,
         \add_0_root_add_0_root_add_446_3/carry[12] ,
         \add_0_root_add_0_root_add_446_3/carry[11] ,
         \add_0_root_add_0_root_add_446_3/carry[10] ,
         \add_0_root_add_0_root_add_446_3/carry[9] ,
         \add_0_root_add_0_root_add_446_3/carry[8] ,
         \add_0_root_add_0_root_add_446_3/carry[7] ,
         \add_0_root_add_0_root_add_446_3/carry[6] ,
         \add_0_root_add_0_root_add_446_3/carry[5] ,
         \add_0_root_add_0_root_add_446_3/carry[4] ,
         \add_0_root_add_0_root_add_446_3/carry[3] , \r1712/carry[3] ,
         \r1712/carry[4] , \add_0_root_add_0_root_add_609_4_cf/carry[19] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[18] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[17] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[16] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[15] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[14] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[13] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[12] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[11] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[10] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[9] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[8] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[7] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[6] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[5] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[4] ,
         \add_0_root_add_0_root_add_609_4_cf/carry[3] , \sub_609/carry[4] ,
         \sub_2_root_sub_0_root_add_266_3/carry[3] ,
         \sub_2_root_sub_0_root_add_266_3/carry[4] ,
         \sub_2_root_sub_0_root_add_266_3/carry[5] ,
         \sub_2_root_sub_0_root_add_266_3/carry[6] ,
         \sub_2_root_sub_0_root_add_266_3/carry[7] ,
         \sub_2_root_sub_0_root_add_266_3/carry[8] ,
         \sub_2_root_sub_0_root_add_266_3/carry[9] , n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3012, n3013,
         n3014, n3015, n3016, n3017, n3019, n3021, n3023, n3025, n3027, n3029,
         n3031, n3033, n3035, n3037, n3039, n3041, n3043, n3045, n3059, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945;
  wire   [15:0] offset_w;
  wire   [19:0] pic_A;
  wire   [2:0] tick;
  wire   [6:0] hour;
  wire   [6:0] min;
  wire   [6:0] sec;
  wire   [2:0] state;
  wire   [2:0] pic_num;
  wire   [9:0] pic_size;
  wire   [19:0] cycle;
  wire   [7:0] count;
  wire   [6:0] hour_n;
  wire   [6:0] min_n;
  wire   [19:0] cycle_n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  DFFRX4 \min_reg[0]  ( .D(min_n[0]), .CK(clk), .RN(n3136), .Q(N6160), .QN(
        n4810) );
  DFFRX4 \min_reg[1]  ( .D(min_n[1]), .CK(clk), .RN(n3125), .Q(N6150), .QN(
        n4869) );
  DFFRX4 \min_reg[4]  ( .D(min_n[4]), .CK(clk), .RN(n3125), .Q(min[4]), .QN(
        n4866) );
  DFFRX1 \tick_reg[0]  ( .D(n1689), .CK(clk), .RN(n3137), .Q(tick[0]) );
  DFFRX1 \tick_reg[1]  ( .D(n1688), .CK(clk), .RN(n3138), .Q(tick[1]), .QN(
        n2980) );
  DFFRX1 \tick_reg[2]  ( .D(n1687), .CK(clk), .RN(n1425), .Q(tick[2]) );
  DFFRX1 \count_reg[0]  ( .D(n1686), .CK(clk), .RN(n3137), .Q(N6482), .QN(
        n1424) );
  DFFRX1 \IM_A_reg[0]  ( .D(n1685), .CK(clk), .RN(n3135), .QN(n1423) );
  DFFRX1 \count_reg[1]  ( .D(n1684), .CK(clk), .RN(n3135), .Q(N6483), .QN(
        n4875) );
  DFFRX1 \IM_A_reg[1]  ( .D(n1683), .CK(clk), .RN(n3140), .QN(n4843) );
  DFFRX1 \count_reg[2]  ( .D(n1682), .CK(clk), .RN(n3135), .Q(N6484), .QN(
        n4874) );
  DFFRX1 \pic_size_reg[7]  ( .D(n1681), .CK(clk), .RN(n3130), .Q(pic_size[7]), 
        .QN(n2965) );
  DFFRX1 \pix_c_reg[0]  ( .D(n1680), .CK(clk), .RN(n3128), .Q(N4429), .QN(
        n4854) );
  DFFRX1 \state_reg[2]  ( .D(n1675), .CK(clk), .RN(n3131), .Q(state[2]), .QN(
        n2963) );
  DFFRX1 flag_512_reg ( .D(n1673), .CK(clk), .RN(n3136), .QN(n1927) );
  DFFRX1 \state_reg[1]  ( .D(n1670), .CK(clk), .RN(n3136), .Q(state[1]), .QN(
        n2957) );
  DFFRX1 \count_reg[3]  ( .D(n1669), .CK(clk), .RN(n3137), .Q(count[3]), .QN(
        n4873) );
  DFFRX1 \count_reg[4]  ( .D(n1668), .CK(clk), .RN(n3135), .Q(count[4]) );
  DFFRX1 \count_reg[5]  ( .D(n1667), .CK(clk), .RN(n3136), .Q(count[5]), .QN(
        n4872) );
  DFFRX1 \count_reg[6]  ( .D(n1666), .CK(clk), .RN(n3138), .Q(count[6]), .QN(
        n4870) );
  DFFRX1 \count_reg[7]  ( .D(n1665), .CK(clk), .RN(n3137), .Q(count[7]), .QN(
        n4871) );
  DFFRX1 \pic_size_reg[9]  ( .D(n1663), .CK(clk), .RN(n3130), .Q(pic_size[9]), 
        .QN(n2958) );
  DFFRX1 \pic_size_reg[8]  ( .D(n1662), .CK(clk), .RN(n3130), .Q(pic_size[8]), 
        .QN(n2974) );
  DFFRX1 \pic_size_reg[6]  ( .D(n1661), .CK(clk), .RN(n3130), .Q(pic_size[6])
         );
  DFFRX1 \pic_size_reg[5]  ( .D(n1660), .CK(clk), .RN(n3131), .Q(pic_size[5])
         );
  DFFRX1 \pic_size_reg[4]  ( .D(n1659), .CK(clk), .RN(n3131), .Q(pic_size[4])
         );
  DFFRX1 \pic_size_reg[3]  ( .D(n1658), .CK(clk), .RN(n3131), .Q(pic_size[3])
         );
  DFFRX1 \pic_size_reg[2]  ( .D(n1657), .CK(clk), .RN(n3131), .Q(pic_size[2]), 
        .QN(n2959) );
  DFFRX1 \pic_size_reg[1]  ( .D(n1656), .CK(clk), .RN(n3131), .Q(pic_size[1]), 
        .QN(n2967) );
  DFFRX1 \pic_size_reg[0]  ( .D(n1655), .CK(clk), .RN(n3131), .Q(N1239), .QN(
        n2975) );
  DFFRX1 flag_128_reg ( .D(n1654), .CK(clk), .RN(n3135), .Q(n2979), .QN(n2016)
         );
  DFFRX1 \offset_reg[0]  ( .D(n1653), .CK(clk), .RN(n3138), .Q(N789), .QN(
        n3082) );
  DFFRX1 \offset_reg[8]  ( .D(n1645), .CK(clk), .RN(n3125), .Q(N797), .QN(
        n3123) );
  DFFRX1 \offset_reg[7]  ( .D(n1644), .CK(clk), .RN(n3135), .Q(N796), .QN(
        n3078) );
  DFFRX1 \offset_reg[6]  ( .D(n1643), .CK(clk), .RN(n3138), .Q(N795), .QN(
        n3076) );
  DFFRX1 \offset_reg[5]  ( .D(n1642), .CK(clk), .RN(n3137), .Q(N794), .QN(
        n3080) );
  DFFRX1 \offset_reg[4]  ( .D(n1641), .CK(clk), .RN(n3135), .Q(N793), .QN(
        n3074) );
  DFFRX1 \offset_reg[2]  ( .D(n1639), .CK(clk), .RN(n3135), .Q(N791), .QN(
        n2968) );
  DFFRX1 \offset_reg[1]  ( .D(n1638), .CK(clk), .RN(n3135), .Q(N790), .QN(
        n2961) );
  DFFRX1 \sec_reg[6]  ( .D(n1619), .CK(clk), .RN(n3141), .Q(sec[6]), .QN(n2978) );
  DFFRX1 \pic_num_reg[2]  ( .D(n1618), .CK(clk), .RN(n3129), .Q(pic_num[2]), 
        .QN(n2984) );
  DFFRX1 \pic_num_reg[1]  ( .D(n1617), .CK(clk), .RN(n3129), .Q(pic_num[1]) );
  DFFRX1 \pic_num_reg[0]  ( .D(n1616), .CK(clk), .RN(n3129), .Q(pic_num[0]), 
        .QN(n2991) );
  DFFRX1 \pic_c_reg[0]  ( .D(n1615), .CK(clk), .RN(n3129), .Q(n4788), .QN(
        n2981) );
  DFFRX1 \pic_c_reg[1]  ( .D(n1614), .CK(clk), .RN(n3129), .Q(n4787), .QN(
        n2983) );
  DFFRX1 \CR_A_reg[0]  ( .D(n1593), .CK(clk), .RN(n3134), .QN(n1420) );
  DFFRX1 \CR_A_reg[1]  ( .D(n1592), .CK(clk), .RN(n3134), .QN(n1419) );
  DFFRX1 \CR_A_reg[2]  ( .D(n1591), .CK(clk), .RN(n3141), .QN(n1418) );
  DFFRX1 \CR_A_reg[3]  ( .D(n1590), .CK(clk), .RN(n3134), .QN(n1417) );
  DFFRX1 \CR_A_reg[4]  ( .D(n1589), .CK(clk), .RN(n3134), .QN(n1416) );
  DFFRX1 \CR_A_reg[5]  ( .D(n1588), .CK(clk), .RN(n3134), .QN(n1415) );
  DFFRX1 \CR_A_reg[6]  ( .D(n1587), .CK(clk), .RN(n3134), .QN(n1414) );
  DFFRX1 \CR_A_reg[7]  ( .D(n1586), .CK(clk), .RN(n3134), .QN(n1413) );
  DFFRX1 \CR_A_reg[8]  ( .D(n1585), .CK(clk), .RN(n3134), .QN(n1412) );
  DFFRX1 \IM_D_t_reg[3][9]  ( .D(n1584), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][9] ), .QN(n2110) );
  DFFRX1 \IM_D_t_reg[3][8]  ( .D(n1583), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][8] ), .QN(n2111) );
  DFFRX1 \IM_D_t_reg[3][7]  ( .D(n1582), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][7] ), .QN(n2112) );
  DFFRX1 \IM_D_t_reg[3][6]  ( .D(n1581), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][6] ), .QN(n2113) );
  DFFRX1 \IM_D_t_reg[3][5]  ( .D(n1580), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][5] ), .QN(n2114) );
  DFFRX1 \IM_D_t_reg[3][4]  ( .D(n1579), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][4] ), .QN(n2115) );
  DFFRX1 \IM_D_t_reg[3][3]  ( .D(n1578), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[3][3] ), .QN(n2116) );
  DFFRX1 \IM_D_t_reg[3][2]  ( .D(n1577), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[3][2] ), .QN(n2117) );
  DFFRX1 \IM_D_t_reg[3][23]  ( .D(n1576), .CK(clk), .RN(n3135), .Q(
        \IM_D_t[3][23] ), .QN(n2118) );
  DFFRX1 \IM_D_t_reg[3][22]  ( .D(n1575), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[3][22] ), .QN(n2119) );
  DFFRX1 \IM_D_t_reg[3][21]  ( .D(n1574), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[3][21] ), .QN(n2120) );
  DFFRX1 \IM_D_t_reg[3][20]  ( .D(n1573), .CK(clk), .RN(n3136), .Q(
        \IM_D_t[3][20] ), .QN(n2121) );
  DFFRX1 \IM_D_t_reg[3][1]  ( .D(n1572), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[3][1] ), .QN(n2122) );
  DFFRX1 \IM_D_t_reg[3][19]  ( .D(n1571), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[3][19] ), .QN(n2123) );
  DFFRX1 \IM_D_t_reg[3][18]  ( .D(n1570), .CK(clk), .RN(n3138), .Q(
        \IM_D_t[3][18] ), .QN(n2124) );
  DFFRX1 \IM_D_t_reg[3][17]  ( .D(n1569), .CK(clk), .RN(n1425), .Q(
        \IM_D_t[3][17] ), .QN(n2125) );
  DFFRX1 \IM_D_t_reg[3][16]  ( .D(n1568), .CK(clk), .RN(n1425), .Q(
        \IM_D_t[3][16] ), .QN(n2126) );
  DFFRX1 \IM_D_t_reg[3][15]  ( .D(n1567), .CK(clk), .RN(n1425), .Q(
        \IM_D_t[3][15] ), .QN(n2127) );
  DFFRX1 \IM_D_t_reg[3][14]  ( .D(n1566), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[3][14] ), .QN(n2128) );
  DFFRX1 \IM_D_t_reg[3][13]  ( .D(n1565), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[3][13] ), .QN(n2129) );
  DFFRX1 \IM_D_t_reg[3][12]  ( .D(n1564), .CK(clk), .RN(n3137), .Q(
        \IM_D_t[3][12] ), .QN(n2130) );
  DFFRX1 \IM_D_t_reg[3][11]  ( .D(n1563), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[3][11] ), .QN(n2131) );
  DFFRX1 \IM_D_t_reg[3][10]  ( .D(n1562), .CK(clk), .RN(n3135), .Q(
        \IM_D_t[3][10] ), .QN(n2132) );
  DFFRX1 \IM_D_t_reg[3][0]  ( .D(n1561), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[3][0] ), .QN(n2133) );
  DFFRX1 \IM_D_t_reg[2][23]  ( .D(n1560), .CK(clk), .RN(n3136), .Q(
        \IM_D_t[2][23] ), .QN(n2068) );
  DFFRX1 \IM_D_t_reg[2][22]  ( .D(n1559), .CK(clk), .RN(n3138), .Q(
        \IM_D_t[2][22] ), .QN(n2069) );
  DFFRX1 \IM_D_t_reg[2][21]  ( .D(n1558), .CK(clk), .RN(n3137), .Q(
        \IM_D_t[2][21] ), .QN(n2070) );
  DFFRX1 \IM_D_t_reg[2][20]  ( .D(n1557), .CK(clk), .RN(n3129), .Q(
        \IM_D_t[2][20] ), .QN(n2071) );
  DFFRX1 \IM_D_t_reg[2][19]  ( .D(n1556), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][19] ), .QN(n2072) );
  DFFRX1 \IM_D_t_reg[2][18]  ( .D(n1555), .CK(clk), .RN(n3131), .Q(
        \IM_D_t[2][18] ), .QN(n2073) );
  DFFRX1 \IM_D_t_reg[2][17]  ( .D(n1554), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][17] ), .QN(n2074) );
  DFFRX1 \IM_D_t_reg[2][16]  ( .D(n1553), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][16] ), .QN(n2075) );
  DFFRX1 \IM_D_t_reg[2][15]  ( .D(n1552), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][15] ), .QN(n2076) );
  DFFRX1 \IM_D_t_reg[2][14]  ( .D(n1551), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][14] ), .QN(n2077) );
  DFFRX1 \IM_D_t_reg[2][13]  ( .D(n1550), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][13] ), .QN(n2078) );
  DFFRX1 \IM_D_t_reg[2][12]  ( .D(n1549), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][12] ), .QN(n2079) );
  DFFRX1 \IM_D_t_reg[2][11]  ( .D(n1548), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][11] ), .QN(n2080) );
  DFFRX1 \IM_D_t_reg[2][10]  ( .D(n1547), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][10] ), .QN(n2081) );
  DFFRX1 \IM_D_t_reg[2][9]  ( .D(n1546), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][9] ), .QN(n2082) );
  DFFRX1 \IM_D_t_reg[2][8]  ( .D(n1545), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][8] ), .QN(n2083) );
  DFFRX1 \IM_D_t_reg[2][7]  ( .D(n1544), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][7] ), .QN(n4746) );
  DFFRX1 \IM_D_t_reg[2][6]  ( .D(n1543), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][6] ), .QN(n4747) );
  DFFRX1 \IM_D_t_reg[2][5]  ( .D(n1542), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][5] ), .QN(n4748) );
  DFFRX1 \IM_D_t_reg[2][4]  ( .D(n1541), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][4] ), .QN(n4749) );
  DFFRX1 \IM_D_t_reg[2][3]  ( .D(n1540), .CK(clk), .RN(n3126), .Q(
        \IM_D_t[2][3] ), .QN(n4750) );
  DFFRX1 \IM_D_t_reg[2][2]  ( .D(n1539), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[2][2] ), .QN(n4751) );
  DFFRX1 \IM_D_t_reg[2][1]  ( .D(n1538), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[2][1] ), .QN(n4752) );
  DFFRX1 \IM_D_t_reg[2][0]  ( .D(n1537), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[2][0] ), .QN(n4753) );
  DFFRX1 \IM_D_t_reg[1][23]  ( .D(n1536), .CK(clk), .RN(n3137), .Q(
        \IM_D_t[1][23] ), .QN(n4762) );
  DFFRX1 \IM_D_t_reg[1][22]  ( .D(n1535), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[1][22] ), .QN(n4763) );
  DFFRX1 \IM_D_t_reg[1][21]  ( .D(n1534), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[1][21] ), .QN(n4764) );
  DFFRX1 \IM_D_t_reg[1][20]  ( .D(n1533), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[1][20] ), .QN(n4765) );
  DFFRX1 \IM_D_t_reg[1][19]  ( .D(n1532), .CK(clk), .RN(n3135), .Q(
        \IM_D_t[1][19] ), .QN(n4767) );
  DFFRX1 \IM_D_t_reg[1][18]  ( .D(n1531), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[1][18] ), .QN(n4768) );
  DFFRX1 \IM_D_t_reg[1][17]  ( .D(n1530), .CK(clk), .RN(n3136), .Q(
        \IM_D_t[1][17] ), .QN(n4769) );
  DFFRX1 \IM_D_t_reg[1][16]  ( .D(n1529), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[1][16] ), .QN(n4770) );
  DFFRX1 \IM_D_t_reg[1][15]  ( .D(n1528), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[1][15] ), .QN(n4771) );
  DFFRX1 \IM_D_t_reg[1][14]  ( .D(n1527), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[1][14] ), .QN(n4772) );
  DFFRX1 \IM_D_t_reg[1][13]  ( .D(n1526), .CK(clk), .RN(n3138), .Q(
        \IM_D_t[1][13] ), .QN(n4773) );
  DFFRX1 \IM_D_t_reg[1][12]  ( .D(n1525), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[1][12] ), .QN(n4774) );
  DFFRX1 \IM_D_t_reg[1][11]  ( .D(n1524), .CK(clk), .RN(n3140), .Q(
        \IM_D_t[1][11] ), .QN(n4775) );
  DFFRX1 \IM_D_t_reg[1][10]  ( .D(n1523), .CK(clk), .RN(n3137), .Q(
        \IM_D_t[1][10] ), .QN(n4776) );
  DFFRX1 \IM_D_t_reg[1][9]  ( .D(n1522), .CK(clk), .RN(n3139), .Q(
        \IM_D_t[1][9] ), .QN(n4754) );
  DFFRX1 \IM_D_t_reg[1][8]  ( .D(n1521), .CK(clk), .RN(n3141), .Q(
        \IM_D_t[1][8] ), .QN(n4755) );
  DFFRX1 \IM_D_t_reg[1][7]  ( .D(n1520), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][7] ), .QN(n4756) );
  DFFRX1 \IM_D_t_reg[1][6]  ( .D(n1519), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][6] ), .QN(n4757) );
  DFFRX1 \IM_D_t_reg[1][5]  ( .D(n1518), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][5] ), .QN(n4758) );
  DFFRX1 \IM_D_t_reg[1][4]  ( .D(n1517), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][4] ), .QN(n4759) );
  DFFRX1 \IM_D_t_reg[1][3]  ( .D(n1516), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][3] ), .QN(n4760) );
  DFFRX1 \IM_D_t_reg[1][2]  ( .D(n1515), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][2] ), .QN(n4761) );
  DFFRX1 \IM_D_t_reg[1][1]  ( .D(n1514), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][1] ), .QN(n4766) );
  DFFRX1 \IM_D_t_reg[1][0]  ( .D(n1513), .CK(clk), .RN(n3133), .Q(
        \IM_D_t[1][0] ), .QN(n4777) );
  DFFRX1 \IM_D_t_reg[0][23]  ( .D(n1512), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][23] ), .QN(n4819) );
  DFFRX1 \IM_D_t_reg[0][22]  ( .D(n1511), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][22] ), .QN(n4820) );
  DFFRX1 \IM_D_t_reg[0][21]  ( .D(n1510), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][21] ), .QN(n4821) );
  DFFRX1 \IM_D_t_reg[0][20]  ( .D(n1509), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][20] ), .QN(n4822) );
  DFFRX1 \IM_D_t_reg[0][19]  ( .D(n1508), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][19] ), .QN(n4824) );
  DFFRX1 \IM_D_t_reg[0][18]  ( .D(n1507), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][18] ), .QN(n4825) );
  DFFRX1 \IM_D_t_reg[0][17]  ( .D(n1506), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][17] ), .QN(n4826) );
  DFFRX1 \IM_D_t_reg[0][16]  ( .D(n1505), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][16] ), .QN(n4827) );
  DFFRX1 \IM_D_t_reg[0][15]  ( .D(n1504), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][15] ), .QN(n4828) );
  DFFRX1 \IM_D_t_reg[0][14]  ( .D(n1503), .CK(clk), .RN(n3127), .Q(
        \IM_D_t[0][14] ), .QN(n4829) );
  DFFRX1 \IM_D_t_reg[0][13]  ( .D(n1502), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][13] ), .QN(n4830) );
  DFFRX1 \IM_D_t_reg[0][12]  ( .D(n1501), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][12] ), .QN(n4831) );
  DFFRX1 \IM_D_t_reg[0][11]  ( .D(n1500), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][11] ), .QN(n4832) );
  DFFRX1 \IM_D_t_reg[0][10]  ( .D(n1499), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][10] ), .QN(n4833) );
  DFFRX1 \IM_D_t_reg[0][9]  ( .D(n1498), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][9] ), .QN(n4811) );
  DFFRX1 \IM_D_t_reg[0][8]  ( .D(n1497), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][8] ), .QN(n4778) );
  DFFRX1 \IM_D_t_reg[0][7]  ( .D(n1496), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][7] ), .QN(n4779) );
  DFFRX1 \IM_D_t_reg[0][6]  ( .D(n1495), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][6] ), .QN(n4780) );
  DFFRX1 \IM_D_t_reg[0][5]  ( .D(n1494), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][5] ), .QN(n4781) );
  DFFRX1 \IM_D_t_reg[0][4]  ( .D(n1493), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][4] ), .QN(n4782) );
  DFFRX1 \IM_D_t_reg[0][3]  ( .D(n1492), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][3] ), .QN(n4783) );
  DFFRX1 \IM_D_t_reg[0][2]  ( .D(n1491), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][2] ), .QN(n4784) );
  DFFRX1 \IM_D_t_reg[0][1]  ( .D(n1490), .CK(clk), .RN(n3129), .Q(
        \IM_D_t[0][1] ), .QN(n4785) );
  DFFRX1 \IM_D_t_reg[0][0]  ( .D(n1489), .CK(clk), .RN(n3128), .Q(
        \IM_D_t[0][0] ), .QN(n4786) );
  DFFRX1 \IM_D_reg[1]  ( .D(n1488), .CK(clk), .RN(n3132), .Q(n4985), .QN(n4823) );
  DFFRX1 \IM_D_reg[2]  ( .D(n1487), .CK(clk), .RN(n3132), .Q(n4984), .QN(n4818) );
  DFFRX1 \IM_D_reg[3]  ( .D(n1486), .CK(clk), .RN(n3132), .Q(n4983), .QN(n4817) );
  DFFRX1 \IM_D_reg[4]  ( .D(n1485), .CK(clk), .RN(n3132), .Q(n4982), .QN(n4816) );
  DFFRX1 \IM_D_reg[5]  ( .D(n1484), .CK(clk), .RN(n3132), .Q(n4981), .QN(n4815) );
  DFFRX1 \IM_D_reg[6]  ( .D(n1483), .CK(clk), .RN(n3132), .Q(n4980), .QN(n4814) );
  DFFRX1 \IM_D_reg[7]  ( .D(n1482), .CK(clk), .RN(n3132), .Q(n4979), .QN(n4813) );
  DFFRX1 \IM_D_reg[8]  ( .D(n1481), .CK(clk), .RN(n3135), .Q(n4978), .QN(n4812) );
  DFFRX1 \IM_D_reg[9]  ( .D(n1480), .CK(clk), .RN(n3132), .Q(n4977), .QN(n3017) );
  DFFRX1 \IM_D_reg[10]  ( .D(n1479), .CK(clk), .RN(n3132), .Q(n4976), .QN(
        n3019) );
  DFFRX1 \IM_D_reg[11]  ( .D(n1478), .CK(clk), .RN(n3132), .Q(n4975), .QN(
        n3021) );
  DFFRX1 \IM_D_reg[12]  ( .D(n1477), .CK(clk), .RN(n3132), .Q(n4974), .QN(
        n3023) );
  DFFRX1 \IM_D_reg[13]  ( .D(n1476), .CK(clk), .RN(n3132), .Q(n4973), .QN(
        n3025) );
  DFFRX1 \IM_D_reg[14]  ( .D(n1475), .CK(clk), .RN(n3132), .Q(n4972), .QN(
        n3027) );
  DFFRX1 \IM_D_reg[15]  ( .D(n1474), .CK(clk), .RN(n3132), .Q(n4971), .QN(
        n3029) );
  DFFRX1 \IM_D_reg[16]  ( .D(n1473), .CK(clk), .RN(n3132), .Q(n4970), .QN(
        n3031) );
  DFFRX1 \IM_D_reg[17]  ( .D(n1472), .CK(clk), .RN(n3132), .Q(n4969), .QN(
        n3033) );
  DFFRX1 \IM_D_reg[18]  ( .D(n1471), .CK(clk), .RN(n3132), .Q(n4968), .QN(
        n3035) );
  DFFRX1 \IM_D_reg[19]  ( .D(n1470), .CK(clk), .RN(n3132), .Q(n4967), .QN(
        n3037) );
  DFFRX1 \IM_D_reg[20]  ( .D(n1469), .CK(clk), .RN(n3134), .Q(n4966), .QN(
        n3039) );
  DFFRX1 \IM_D_reg[21]  ( .D(n1468), .CK(clk), .RN(n3134), .Q(n4965), .QN(
        n3041) );
  DFFRX1 \IM_D_reg[22]  ( .D(n1467), .CK(clk), .RN(n3134), .Q(n4964), .QN(
        n3043) );
  DFFRX1 \IM_D_reg[23]  ( .D(n1466), .CK(clk), .RN(n3134), .Q(n4963), .QN(
        n3045) );
  DFFRX1 \IM_D_reg[0]  ( .D(n1465), .CK(clk), .RN(n3134), .Q(n4986), .QN(n4834) );
  DFFSX1 IM_WEN_reg ( .D(n1464), .CK(clk), .SN(n3133), .QN(n2098) );
  DFFRX1 \pic_A_reg[19]  ( .D(n1463), .CK(clk), .RN(n3131), .Q(pic_A[19]), 
        .QN(n4717) );
  DFFRX1 \pic_A_reg[4]  ( .D(n1448), .CK(clk), .RN(n3129), .Q(pic_A[4]), .QN(
        n4713) );
  DFFRX1 \pic_A_reg[3]  ( .D(n1447), .CK(clk), .RN(n3128), .Q(pic_A[3]), .QN(
        n4714) );
  DFFRX1 \pic_A_reg[2]  ( .D(n1446), .CK(clk), .RN(n3128), .Q(pic_A[2]), .QN(
        n4715) );
  DFFRX1 \IM_A_reg[3]  ( .D(n1443), .CK(clk), .RN(n3141), .QN(n4841) );
  DFFRX1 \IM_A_reg[4]  ( .D(n1442), .CK(clk), .RN(n3141), .QN(n4840) );
  DFFRX1 \IM_A_reg[5]  ( .D(n1441), .CK(clk), .RN(n3141), .QN(n4839) );
  DFFRX1 \IM_A_reg[6]  ( .D(n1440), .CK(clk), .RN(n3141), .QN(n4838) );
  DFFRX1 \IM_A_reg[7]  ( .D(n1439), .CK(clk), .RN(n3141), .QN(n4837) );
  DFFRX1 \IM_A_reg[8]  ( .D(n1438), .CK(clk), .RN(n3138), .Q(n4962), .QN(n4836) );
  DFFRX1 \IM_A_reg[9]  ( .D(n1437), .CK(clk), .RN(n3141), .Q(n4961), .QN(n4835) );
  DFFRX1 \IM_A_reg[10]  ( .D(n1436), .CK(clk), .RN(n3139), .Q(n4960), .QN(
        n4853) );
  DFFRX1 \IM_A_reg[11]  ( .D(n1435), .CK(clk), .RN(n3140), .Q(n4959), .QN(
        n4852) );
  DFFRX1 \IM_A_reg[12]  ( .D(n1434), .CK(clk), .RN(n3139), .Q(n4958), .QN(
        n4851) );
  DFFRX1 \IM_A_reg[13]  ( .D(n1433), .CK(clk), .RN(n3140), .Q(n4957), .QN(
        n4850) );
  DFFRX1 \IM_A_reg[14]  ( .D(n1432), .CK(clk), .RN(n1425), .Q(n4956), .QN(
        n4849) );
  DFFRX1 \IM_A_reg[15]  ( .D(n1431), .CK(clk), .RN(n3139), .Q(n4955), .QN(
        n4848) );
  DFFRX1 \IM_A_reg[16]  ( .D(n1430), .CK(clk), .RN(n3127), .Q(n4954), .QN(
        n4847) );
  DFFRX1 \IM_A_reg[17]  ( .D(n1429), .CK(clk), .RN(n3140), .Q(n4953), .QN(
        n4846) );
  DFFRX1 \IM_A_reg[18]  ( .D(n1428), .CK(clk), .RN(n3139), .Q(n4952), .QN(
        n4845) );
  DFFRX1 \IM_A_reg[19]  ( .D(n1427), .CK(clk), .RN(n3131), .Q(n4951), .QN(
        n4844) );
  DFFRX1 \IM_A_reg[2]  ( .D(n1426), .CK(clk), .RN(n3141), .QN(n4842) );
  DPA_DW01_add_0 add_0_root_add_536_3_cf ( .A({1'b0, 1'b0, 1'b0, 
        offset_w[15:8], N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, 
        1'b0}), .B({N7645, N7646, N7647, N7648, N7649, N7650, N7651, N7652, 
        N7653, N7654, N7655, N7656, N7657, N7658, N7659, N7660, N7661, N7662, 
        N7663, N7664}), .CI(1'b0), .SUM({N3771, N3770, N3769, N3768, N3767, 
        N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, 
        N3756, N3755, N3754, N3753, N3752}) );
  DPA_DW01_add_1 add_0_root_add_519_3_cf ( .A({1'b0, 1'b0, 1'b0, 
        offset_w[15:8], N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, 
        1'b0}), .B({N7625, N7626, N7627, N7628, N7629, N7630, N7631, N7632, 
        N7633, N7634, N7635, N7636, N7637, N7638, N7639, N7640, N7641, N7642, 
        N7643, N7644}), .CI(1'b0), .SUM({N3636, N3635, N3634, N3633, N3632, 
        N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, 
        N3621, N3620, N3619, N3618, N3617}) );
  DPA_DW01_inc_0 add_993 ( .A({hour[6:2], N5926, N5910}), .SUM({N6810, N6809, 
        N6808, N6807, N6806, N6805, N6804}) );
  DPA_DW01_inc_1 add_989 ( .A({min[6:3], N6151, N6150, N6160}), .SUM({N6789, 
        N6788, N6787, N6786, N6785, N6784, N6783}) );
  DPA_DW01_inc_2 add_984 ( .A({sec[6:3], N6392, N6391, N6401}), .SUM({N6775, 
        N6774, N6773, N6772, N6771, N6770, N6769}) );
  DPA_DW01_inc_3 add_980 ( .A(cycle), .SUM({N6764, N6763, N6762, N6761, N6760, 
        N6759, N6758, N6757, N6756, N6755, N6754, N6753, N6752, N6751, N6750, 
        N6749, N6748, N6747, N6746, N6745}) );
  DPA_DW01_add_3 add_0_root_add_656_2 ( .A({1'b0, 1'b0, N804, N803, N802, N801, 
        N800, N799, N798, n3073, n3079, n3077, N794, n3075, n3016, n3071, 
        n3072, n3083, 1'b0, 1'b0}), .B({N4105, N4104, N4103, N4102, N4101, 
        N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, 
        N4090, N4089, N4088, N4087, N4086}), .CI(1'b0), .SUM({N4995, N4994, 
        N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, 
        N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976}) );
  DPA_DW01_add_4 add_634 ( .A({offset_w[15:8], N4352, N4351, N4350, N4349, 
        N4348, N4347, N4346, N4345}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .CI(1'b0), .SUM({N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, 
        N4636, N4635, N4634, N4633, N4632, N4631}) );
  DPA_DW01_add_5 add_633 ( .A({N804, N803, N802, N801, N800, N799, N798, n3073, 
        n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0}), .CI(1'b0), .SUM({N4630, N4629, N4628, N4627, N4626, 
        N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, 
        N4615}) );
  DPA_DW01_add_6 add_594 ( .A({1'b0, \IM_D_t[1][23] , \IM_D_t[1][22] , 
        \IM_D_t[1][21] , \IM_D_t[1][20] , \IM_D_t[1][19] , \IM_D_t[1][18] , 
        \IM_D_t[1][17] , \IM_D_t[1][16] , \IM_D_t[1][15] , \IM_D_t[1][14] , 
        \IM_D_t[1][13] , \IM_D_t[1][12] , \IM_D_t[1][11] , \IM_D_t[1][10] , 
        \IM_D_t[1][9] , \IM_D_t[1][8] , \IM_D_t[1][7] , \IM_D_t[1][6] , 
        \IM_D_t[1][5] , \IM_D_t[1][4] , \IM_D_t[1][3] , \IM_D_t[1][2] , 
        \IM_D_t[1][1] , \IM_D_t[1][0] }), .B({1'b0, \IM_D_t[3][23] , 
        \IM_D_t[3][22] , \IM_D_t[3][21] , \IM_D_t[3][20] , \IM_D_t[3][19] , 
        \IM_D_t[3][18] , \IM_D_t[3][17] , \IM_D_t[3][16] , \IM_D_t[3][15] , 
        \IM_D_t[3][14] , \IM_D_t[3][13] , \IM_D_t[3][12] , \IM_D_t[3][11] , 
        \IM_D_t[3][10] , \IM_D_t[3][9] , \IM_D_t[3][8] , \IM_D_t[3][7] , 
        \IM_D_t[3][6] , \IM_D_t[3][5] , \IM_D_t[3][4] , \IM_D_t[3][3] , 
        \IM_D_t[3][2] , \IM_D_t[3][1] , \IM_D_t[3][0] }), .CI(1'b0), .SUM({
        N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, 
        N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, 
        N4274, N4273, N4272, N4271, SYNOPSYS_UNCONNECTED__0}) );
  DPA_DW01_add_7 add_0_root_add_571_2 ( .A({1'b0, 1'b0, 1'b0, offset_w[15:8], 
        N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, 1'b0}), .B({
        N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, 
        N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086}), 
        .CI(1'b0), .SUM({N4125, N4124, N4123, N4122, N4121, N4120, N4119, 
        N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, 
        N4108, N4107, N4106}) );
  DPA_DW01_sub_0 sub_413 ( .A({N804, N803, N802, N801, N800, N799, N798, n3073, 
        n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .CI(1'b0), .DIFF({N2503, N2502, N2501, N2500, 
        N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, 
        N2489, N2488}) );
  DPA_DW01_sub_1 sub_0_root_sub_192 ( .A({N527, N526, N525, N524, N523, N522, 
        N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, 
        N509, N508}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, pic_size[9:1], N1239}), .CI(1'b0), .DIFF({N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, 
        N551, N550, N549, N548}) );
  DPA_DW01_add_14 r1772 ( .A({1'b0, N4428, N4427, N4426, N4425, N4424, N4423, 
        N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, 
        N4412, N4411, N4410, N4409}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .CI(1'b0), .SUM({N5167, N5166, N5165, N5164, N5163, 
        N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, 
        N5152, N5151, N5150, N5149, N5148, N5147}) );
  DPA_DW01_add_15 r1758 ( .A({N4428, N4427, N4426, N4425, N4424, N4423, N4422, 
        N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, 
        N4411, N4410, N4409}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \gt_332/n9 , 
        \gt_332/n15 , n3305, n3015, 1'b0}), .CI(1'b0), .SUM({N4105, N4104, 
        N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, 
        N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086}) );
  DPA_DW01_add_16 r1756 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .B({N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, 
        N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409}), 
        .CI(1'b0), .SUM({N7645, N7646, N7647, N7648, N7649, N7650, N7651, 
        N7652, N7653, N7654, N7655, N7656, N7657, N7658, N7659, N7660, N7661, 
        N7662, N7663, N7664}) );
  DPA_DW01_add_17 r1753 ( .A({1'b0, 1'b0, \IM_D_t[2][23] , \IM_D_t[2][22] , 
        \IM_D_t[2][21] , \IM_D_t[2][20] , \IM_D_t[2][19] , \IM_D_t[2][18] , 
        \IM_D_t[2][17] , \IM_D_t[2][16] , \IM_D_t[2][15] , \IM_D_t[2][14] , 
        \IM_D_t[2][13] , \IM_D_t[2][12] , \IM_D_t[2][11] , \IM_D_t[2][10] , 
        \IM_D_t[2][9] , \IM_D_t[2][8] , \IM_D_t[2][7] , \IM_D_t[2][6] , 
        \IM_D_t[2][5] , \IM_D_t[2][4] , \IM_D_t[2][3] , \IM_D_t[2][2] , 
        \IM_D_t[2][1] , \IM_D_t[2][0] }), .B({1'b0, 1'b0, \IM_D_t[3][23] , 
        \IM_D_t[3][22] , \IM_D_t[3][21] , \IM_D_t[3][20] , \IM_D_t[3][19] , 
        \IM_D_t[3][18] , \IM_D_t[3][17] , \IM_D_t[3][16] , \IM_D_t[3][15] , 
        \IM_D_t[3][14] , \IM_D_t[3][13] , \IM_D_t[3][12] , \IM_D_t[3][11] , 
        \IM_D_t[3][10] , \IM_D_t[3][9] , \IM_D_t[3][8] , \IM_D_t[3][7] , 
        \IM_D_t[3][6] , \IM_D_t[3][5] , \IM_D_t[3][4] , \IM_D_t[3][3] , 
        \IM_D_t[3][2] , \IM_D_t[3][1] , \IM_D_t[3][0] }), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, N3686, N3685, N3684, N3683, N3682, N3681, 
        N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, 
        N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662}) );
  DPA_DW01_add_18 r1751 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .B({N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, 
        N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409}), 
        .CI(1'b0), .SUM({N7625, N7626, N7627, N7628, N7629, N7630, N7631, 
        N7632, N7633, N7634, N7635, N7636, N7637, N7638, N7639, N7640, N7641, 
        N7642, N7643, N7644}) );
  DPA_DW01_add_19 r1748 ( .A({N804, N803, N802, N801, N800, N799, N798, n3073, 
        n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1}), .CI(1'b0), .SUM({N3228, N3227, N3226, N3225, N3224, 
        N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, 
        N3213}) );
  DPA_DW01_add_20 r1743 ( .A({1'b0, N4428, N4427, N4426, N4425, N4424, N4423, 
        N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, 
        N4412, N4411, N4410, N4409}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b0}), .CI(1'b0), .SUM({N3004, N3003, N3002, N3001, N3000, 
        N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, 
        N2989, N2988, N2987, N2986, N2985, N2984}) );
  DPA_DW01_add_21 r1742 ( .A({N804, N803, N802, N801, N800, N799, N798, n3073, 
        n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1}), .CI(1'b0), .SUM({N2959, N2958, N2957, N2956, N2955, 
        N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, 
        N2944}) );
  DPA_DW01_add_22 r1735 ( .A({N4428, N4427, N4426, N4425, N4424, N4423, N4422, 
        N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, 
        N4411, N4410, N4409}), .B({1'b0, 1'b0, 1'b0, offset_w[15:8], N4352, 
        N4351, N4350, N4349, N4348, N4347, N4346, N4345, 1'b0}), .CI(1'b0), 
        .SUM({N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, 
        N2414, N2413, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, 
        N3732}) );
  DPA_DW01_inc_4 r1734 ( .A({offset_w[15:8], N4352, N4351, N4350, N4349, N4348, 
        N4347, N4346, N4345}), .SUM({n71, n72, n73, n74, n75, n76, n77, n78, 
        n79, n80, n81, n82, n83, n84, n85, n86}) );
  DPA_DW01_inc_5 r1733 ( .A({N804, N803, N802, N801, N800, N799, N798, n3073, 
        n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083}), .SUM({n87, 
        n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
        n102}) );
  DPA_DW01_add_23 r1732 ( .A({1'b0, \IM_D_t[0][23] , \IM_D_t[0][22] , 
        \IM_D_t[0][21] , \IM_D_t[0][20] , \IM_D_t[0][19] , \IM_D_t[0][18] , 
        \IM_D_t[0][17] , \IM_D_t[0][16] , \IM_D_t[0][15] , \IM_D_t[0][14] , 
        \IM_D_t[0][13] , \IM_D_t[0][12] , \IM_D_t[0][11] , \IM_D_t[0][10] , 
        \IM_D_t[0][9] , \IM_D_t[0][8] , \IM_D_t[0][7] , \IM_D_t[0][6] , 
        \IM_D_t[0][5] , \IM_D_t[0][4] , \IM_D_t[0][3] , \IM_D_t[0][2] , 
        \IM_D_t[0][1] , \IM_D_t[0][0] }), .B({1'b0, IM_Q}), .CI(1'b0), .SUM({
        N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, 
        N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, 
        N2185, N2184, N2183, N2182, SYNOPSYS_UNCONNECTED__2}) );
  DPA_DW01_add_24 r1731 ( .A({N4428, N4427, N4426, N4425, N4424, N4423, N4422, 
        N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, 
        N4411, N4410, N4409}), .B({1'b0, 1'b0, 1'b0, offset_w[15:8], N4352, 
        N4351, N4350, N4349, N4348, N4347, N4346, N4345, 1'b0}), .CI(1'b1), 
        .SUM({N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, 
        N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, 
        N2318}) );
  DPA_DW01_sub_2 r1720 ( .A({N886, N885, N884, N883, N882, N881, N880, N879, 
        N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .CI(1'b0), .DIFF({
        N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, 
        N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024})
         );
  DPA_DW01_add_25 r1719 ( .A({1'b0, 1'b0, N804, N803, N802, N801, N800, N799, 
        N798, n3073, n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083, 
        1'b0, 1'b0}), .B({N486, N485, N484, N483, N482, N481, N480, N479, N478, 
        N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467}), 
        .CI(1'b0), .SUM({N963, N962, N961, N960, N959, N958, N957, N956, N955, 
        N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944}) );
  DPA_DW01_add_26 r1718 ( .A({N486, N485, N484, N483, N482, N481, N480, N479, 
        N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467}), .B({1'b0, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, 
        N696, N695, N694, N693, N692, N691, N690, N689}), .CI(1'b0), .SUM({
        N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, 
        N874, N873, N872, N871, N870, N869, N868, N867}) );
  DPA_DW01_add_27 r1714 ( .A({1'b0, 1'b0, N804, N803, N802, N801, N800, N799, 
        N798, n3073, n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083, 
        1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, pic_size[9:1], N1239}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__3, 
        N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, 
        N695, N694, N693, N692, N691, N690, N689}) );
  DPA_DW01_add_28 r1707 ( .A(pic_A), .B({1'b0, 1'b0, 1'b0, 1'b0, N804, N803, 
        N802, N801, N800, N799, N798, n3073, n3079, n3077, n3081, n3075, n3016, 
        n3071, n3072, n3083}), .CI(1'b0), .SUM({N527, N526, N525, N524, N523, 
        N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, 
        N510, N509, N508}) );
  DPA_DW01_add_29 r1706 ( .A({1'b0, 1'b0, 1'b0, 1'b0, N804, N803, N802, N801, 
        N800, N799, N798, n3073, n3079, n3077, n3081, n3075, n3016, n3071, 
        n3072, n3083}), .B({N486, N485, N484, N483, N482, N481, N480, N479, 
        N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467}), .CI(1'b0), .SUM({N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, 
        N496, N495, N494, N493, N492, N491, N490, N489, N488, N487}) );
  DPA_DW01_add_30 r1705 ( .A(pic_A), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \gt_332/n9 , \gt_332/n15 , n3305, n3015}), .CI(1'b0), .SUM({N486, N485, 
        N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, 
        N472, N471, N470, N469, N468, N467}) );
  DPA_DW01_inc_6 r1701 ( .A({count[7:3], N6484, N6483, N6482}), .SUM({n137, 
        n138, n139, n140, n141, n142, n143, n144}) );
  DPA_DW01_add_80 add_1_root_r1754 ( .A({1'b0, 1'b0, \IM_D_t[0][23] , 
        \IM_D_t[0][22] , \IM_D_t[0][21] , \IM_D_t[0][20] , \IM_D_t[0][19] , 
        \IM_D_t[0][18] , \IM_D_t[0][17] , \IM_D_t[0][16] , \IM_D_t[0][15] , 
        \IM_D_t[0][14] , \IM_D_t[0][13] , \IM_D_t[0][12] , \IM_D_t[0][11] , 
        \IM_D_t[0][10] , \IM_D_t[0][9] , \IM_D_t[0][8] , \IM_D_t[0][7] , 
        \IM_D_t[0][6] , \IM_D_t[0][5] , \IM_D_t[0][4] , \IM_D_t[0][3] , 
        \IM_D_t[0][2] , \IM_D_t[0][1] , \IM_D_t[0][0] }), .B({1'b0, 1'b0, 
        \IM_D_t[1][23] , \IM_D_t[1][22] , \IM_D_t[1][21] , \IM_D_t[1][20] , 
        \IM_D_t[1][19] , \IM_D_t[1][18] , \IM_D_t[1][17] , \IM_D_t[1][16] , 
        \IM_D_t[1][15] , \IM_D_t[1][14] , \IM_D_t[1][13] , \IM_D_t[1][12] , 
        \IM_D_t[1][11] , \IM_D_t[1][10] , \IM_D_t[1][9] , \IM_D_t[1][8] , 
        \IM_D_t[1][7] , \IM_D_t[1][6] , \IM_D_t[1][5] , \IM_D_t[1][4] , 
        \IM_D_t[1][3] , \IM_D_t[1][2] , \IM_D_t[1][1] , \IM_D_t[1][0] }), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__4, n4945, n4944, n4943, n4942, 
        n4941, n4940, n4939, n4938, n4937, n4936, n4935, n4934, n4933, n4932, 
        n4931, n4930, n4929, n4928, n4927, n4926, n4925, n4924, n4923, n4922, 
        n4921}) );
  DPA_DW01_add_79 add_0_root_r1754 ( .A({1'b0, N3686, N3685, N3684, N3683, 
        N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, 
        N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, 
        N3662}), .B({1'b0, n4945, n4944, n4943, n4942, n4941, n4940, n4939, 
        n4938, n4937, n4936, n4935, n4934, n4933, n4932, n4931, n4930, n4929, 
        n4928, n4927, n4926, n4925, n4924, n4923, n4922, n4921}), .CI(1'b0), 
        .SUM({N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, 
        N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, 
        N3692, N3691, N3690, N3689, N3688, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  DPA_DW01_add_72 add_2_root_add_0_root_add_446_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({N4428, N4427, N4426, N4425, N4424, N4423, 
        N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, 
        N4412, N4411, N4410, N4409}), .CI(1'b0), .SUM({N2849, N2848, N2847, 
        N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, 
        N2836, N2835, N2834, N2833, N2832, N2831, N2830}) );
  DPA_DW01_add_71 add_1_root_add_0_root_add_446_3 ( .A({N2849, N2848, N2847, 
        N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, 
        N2836, N2835, N2834, N2833, N2832, N2831, N2830}), .B({1'b0, 1'b0, 
        N804, N803, N802, N801, N800, N799, N798, n3073, N796, N795, N794, 
        N793, n3016, n3071, n3072, N789, 1'b0, 1'b0}), .CI(1'b0), .SUM({N2829, 
        N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, 
        N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2850}) );
  DPA_DW01_add_70 add_1_root_add_0_root_add_209_3 ( .A(pic_A), .B({1'b0, N707, 
        N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, 
        N694, N693, N692, N691, N690, N689}), .CI(1'b0), .SUM({N688, N687, 
        N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, 
        N674, N673, N672, N671, N670, N709}) );
  DPA_DW01_add_67 add_1_root_add_0_root_add_661_4_cf ( .A({N7625, N7626, N7627, 
        N7628, N7629, N7630, N7631, N7632, N7633, N7634, N7635, N7636, N7637, 
        N7638, N7639, N7640, N7641, N7642, N7643, N7644}), .B({1'b0, 1'b0, 
        N804, N803, N802, N801, N800, N799, N798, n3073, N796, N795, N794, 
        N793, n3016, n3071, n3072, N789, 1'b0, 1'b0}), .CI(1'b0), .SUM({N7604, 
        N7605, N7606, N7607, N7608, N7609, N7610, N7611, N7612, N7613, N7614, 
        N7615, N7616, N7617, N7618, N7619, N7620, N7621, N7622, N5021}) );
  DPA_DW01_add_66 add_1_root_add_1_root_add_282_4 ( .A(pic_A), .B({1'b0, N707, 
        N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, 
        N694, N693, N692, N691, N690, N689}), .CI(1'b1), .SUM({N1400, N1399, 
        N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, 
        N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1441}) );
  DPA_DW01_add_63 add_1_root_add_0_root_add_579_4_cf ( .A({1'b0, 1'b0, 1'b0, 
        offset_w[15:8], N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, 
        1'b0}), .B({N7625, N7626, N7627, N7628, N7629, N7630, N7631, N7632, 
        N7633, N7634, N7635, N7636, N7637, N7638, N7639, N7640, N7641, N7642, 
        N7643, N7644}), .CI(1'b0), .SUM({N7666, N7667, N7668, N7669, N7670, 
        N7671, N7672, N7673, N7674, N7675, N7676, N7677, N7678, N7679, N7680, 
        N7681, N7682, N7683, N7684, N4176}) );
  DPA_DW01_add_41 add_1_root_add_0_root_add_601_3 ( .A({N4428, N4427, N4426, 
        N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, 
        N4415, N4414, N4413, N4412, N4411, N4410, N4409}), .B({1'b0, 1'b0, 
        n2976, N4360, N4359, N4358, N4357, N4356, N4355, N4354, n4729, N4352, 
        N4351, N4350, N4349, N4348, N4347, N4346, N4345, 1'b0}), .CI(1'b0), 
        .SUM({N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, 
        N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, 
        N4364}) );
  DPA_DW01_add_74 add_1_root_add_0_root_add_609_4_cf ( .A({1'b0, 1'b0, 1'b0, 
        offset_w[15:8], N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, 
        1'b0}), .B({N7645, N7646, N7647, N7648, N7649, N7650, N7651, N7652, 
        N7653, N7654, N7655, N7656, N7657, N7658, N7659, N7660, N7661, N7662, 
        N7663, N7664}), .CI(1'b0), .SUM({N7686, N7687, N7688, N7689, N7690, 
        N7691, N7692, N7693, N7694, N7695, N7696, N7697, N7698, N7699, N7700, 
        N7701, N7702, N7703, N7704, N4454}) );
  DPA_DW01_add_78 add_1_root_sub_0_root_add_266_3 ( .A({n2956, n2956, n2956, 
        n2956, n2956, n2956, n2956, n2956, n2956, n2956, N1248, N1247, N1246, 
        N1245, N1244, N1243, N1242, N1241, n2967, N1239}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N804, N803, N802, N801, N800, N799, N798, n3073, n3079, 
        n3077, n3081, n3075, n3016, n3071, n3072, n3083}), .CI(1'b0), .SUM({
        N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, 
        N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259})
         );
  DPA_DW01_add_77 add_0_root_sub_0_root_add_266_3 ( .A({N1278, N1277, N1276, 
        N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261, N1260, N1259}), .B({N486, N485, 
        N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, 
        N472, N471, N470, N469, N468, N467}), .CI(1'b0), .SUM({N1298, N1297, 
        N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, 
        N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279}) );
  DPA_DW01_add_75 add_0_root_r1717 ( .A({1'b0, 1'b0, N804, N803, N802, N801, 
        N800, N799, N798, n3073, n3079, n3077, n3081, n3075, n3016, n3071, 
        n3072, n3083, 1'b1, 1'b0}), .B({N486, N485, N484, N483, N482, N481, 
        N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, 
        N468, N467}), .CI(1'b0), .SUM({N826, N825, N824, N823, N822, N821, 
        N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, 
        N808, N807}) );
  DPA_DW01_add_44 add_1_root_add_0_root_add_278_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \gt_332/n9 , \gt_332/n15 , n3305, n3015, 1'b0}), .B(pic_A), .CI(1'b0), 
        .SUM({N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, 
        N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, 
        N1336}) );
  DPA_DW01_add_43 add_0_root_add_0_root_add_278_2 ( .A({1'b0, 1'b0, N804, N803, 
        N802, N801, N800, N799, N798, n3073, n3079, n3077, n3081, n3075, n3016, 
        n3071, n3072, n3083, 1'b0, 1'b0}), .B({N1355, N1354, N1353, N1352, 
        N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, 
        N1341, N1340, N1339, N1338, N1337, N1336}), .CI(1'b0), .SUM({N1375, 
        N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, 
        N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356}) );
  DPA_DW01_add_33 add_1_root_r1747 ( .A({1'b0, 1'b0, IM_Q[7:0]}), .B({1'b0, 
        1'b0, \IM_D_t[1][7] , \IM_D_t[1][6] , \IM_D_t[1][5] , \IM_D_t[1][4] , 
        \IM_D_t[1][3] , \IM_D_t[1][2] , \IM_D_t[1][1] , \IM_D_t[1][0] }), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__7, n4898, n4897, n4896, n4895, 
        n4894, n4893, n4892, n4891, n4890}) );
  DPA_DW01_add_32 add_2_root_r1747 ( .A({1'b0, 1'b0, \IM_D_t[2][7] , 
        \IM_D_t[2][6] , \IM_D_t[2][5] , \IM_D_t[2][4] , \IM_D_t[2][3] , 
        \IM_D_t[2][2] , \IM_D_t[2][1] , \IM_D_t[2][0] }), .B({1'b0, 1'b0, 
        \IM_D_t[0][7] , \IM_D_t[0][6] , \IM_D_t[0][5] , \IM_D_t[0][4] , 
        \IM_D_t[0][3] , \IM_D_t[0][2] , \IM_D_t[0][1] , \IM_D_t[0][0] }), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__8, N3162, N3161, N3160, N3159, 
        N3158, N3157, N3156, N3155, N3154}) );
  DPA_DW01_add_31 add_0_root_r1747 ( .A({1'b0, 1'b0, N3162, N3161, N3160, 
        N3159, N3158, N3157, N3156, N3155, N3154}), .B({1'b0, 1'b0, n4898, 
        n4897, n4896, n4895, n4894, n4893, n4892, n4891, n4890}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__9, N3171, N3170, N3169, N3168, N3167, 
        N3166, N3165, N3164, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11}) );
  DPA_DW01_add_46 add_1_root_add_1_root_add_205_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \gt_332/n9 , \gt_332/n15 , n3305, n3015, 1'b0}), .B(pic_A), .CI(1'b1), 
        .SUM({N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, 
        N612, N611, N610, N609, N608, N607, N606, N605, N604}) );
  DPA_DW01_add_45 add_0_root_add_1_root_add_205_3 ( .A({1'b0, 1'b0, N804, N803, 
        N802, N801, N800, N799, N798, n3073, n3079, n3077, n3081, n3075, n3016, 
        n3071, n3072, n3083, 1'b0, 1'b0}), .B({N623, N622, N621, N620, N619, 
        N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, 
        N606, N605, N604}), .CI(1'b0), .SUM({N663, N662, N661, N660, N659, 
        N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, 
        N646, N645, N644}) );
  DPA_DW01_add_48 add_1_root_add_1_root_add_441_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \gt_332/n9 , \gt_332/n15 , n3305, n3015, 1'b0}), .B({N4428, N4427, 
        N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, 
        N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409}), .CI(1'b1), 
        .SUM({N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, 
        N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, 
        N2745}) );
  DPA_DW01_add_47 add_0_root_add_1_root_add_441_3 ( .A({1'b0, 1'b0, N804, N803, 
        N802, N801, N800, N799, N798, n3073, N796, N795, N794, N793, n3016, 
        n3071, n3072, n3083, 1'b0, 1'b0}), .B({N2764, N2763, N2762, N2761, 
        N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, 
        N2750, N2749, N2748, N2747, N2746, N2745}), .CI(1'b0), .SUM({N2804, 
        N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, 
        N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785}) );
  DPA_DW01_add_51 add_2_root_add_0_root_add_869_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N6509, N6508, N6507, 
        N6506, N6505, N6504, n3305, n3015}), .B({N4428, N4427, N4426, N4425, 
        N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, 
        N4414, N4413, N4412, N4411, N4410, N4409}), .CI(1'b0), .SUM({N6549, 
        N6548, N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, 
        N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530}) );
  DPA_DW01_add_50 add_1_root_add_0_root_add_869_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, N6490, N6489, N6488, N6487, 
        N6486, n4873, N6484, N6483, N6482}), .B({N800, N799, N798, n3073, 
        n3079, n3077, n3081, n3075, n3016, n3071, n3072, n3083, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N6529, N6528, 
        N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, 
        N6517, N6516, N6515, N6514, N6513, N6512, N6511, N6510}) );
  DPA_DW01_add_49 add_0_root_add_0_root_add_869_4 ( .A({N6529, N6528, N6527, 
        N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, N6517, 
        N6516, N6515, N6514, N6513, N6512, N6511, N6510}), .B({N6549, N6548, 
        N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, N6538, 
        N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530}), .CI(1'b0), 
        .SUM({N6569, N6568, N6567, N6566, N6565, N6564, N6563, N6562, N6561, 
        N6560, N6559, N6558, N6557, N6556, N6555, N6554, N6553, N6552, N6551, 
        N6550}) );
  ADDHXL \mult_817/U6  ( .A(N6401), .B(N6391), .CO(\mult_817/n5 ), .S(N6294)
         );
  ADDFXL \mult_817/U5  ( .A(N6392), .B(N6391), .CI(\mult_817/n5 ), .CO(
        \mult_817/n4 ), .S(N6295) );
  ADDFXL \mult_817/U4  ( .A(sec[3]), .B(N6392), .CI(\mult_817/n4 ), .CO(
        \mult_817/n3 ), .S(N6296) );
  ADDFXL \mult_817/U3  ( .A(sec[4]), .B(sec[3]), .CI(\mult_817/n3 ), .CO(
        \mult_817/n2 ), .S(N6297) );
  ADDHXL \mult_819/U6  ( .A(N6401), .B(n2994), .CO(\mult_819/n5 ), .S(N6321)
         );
  ADDFXL \mult_819/U5  ( .A(N6311), .B(n2994), .CI(\mult_819/n5 ), .CO(
        \mult_819/n4 ), .S(N6322) );
  ADDFXL \mult_819/U4  ( .A(N6312), .B(N6311), .CI(\mult_819/n4 ), .CO(
        \mult_819/n3 ), .S(N6323) );
  ADDFXL \mult_819/U3  ( .A(N6313), .B(N6312), .CI(\mult_819/n3 ), .CO(
        \mult_819/n2 ), .S(N6324) );
  ADDHXL \mult_821/U6  ( .A(N6401), .B(N6391), .CO(\mult_821/n5 ), .S(N6348)
         );
  ADDFXL \mult_821/U5  ( .A(n2995), .B(N6391), .CI(\mult_821/n5 ), .CO(
        \mult_821/n4 ), .S(N6349) );
  ADDFXL \mult_821/U4  ( .A(N6339), .B(n2995), .CI(\mult_821/n4 ), .CO(
        \mult_821/n3 ), .S(N6350) );
  ADDFXL \mult_821/U3  ( .A(N6340), .B(N6339), .CI(\mult_821/n3 ), .CO(
        \mult_821/n2 ), .S(N6351) );
  ADDHXL \mult_823/U6  ( .A(N6401), .B(n2994), .CO(\mult_823/n5 ), .S(N6375)
         );
  ADDFXL \mult_823/U5  ( .A(N6365), .B(n2994), .CI(\mult_823/n5 ), .CO(
        \mult_823/n4 ), .S(N6376) );
  ADDFXL \mult_823/U4  ( .A(N6366), .B(N6365), .CI(\mult_823/n4 ), .CO(
        \mult_823/n3 ), .S(N6377) );
  ADDFXL \mult_823/U3  ( .A(N6367), .B(N6366), .CI(\mult_823/n3 ), .CO(
        \mult_823/n2 ), .S(N6378) );
  ADDHXL \mult_827/U6  ( .A(N6401), .B(n2994), .CO(\mult_827/n5 ), .S(N6428)
         );
  ADDFXL \mult_827/U5  ( .A(N6418), .B(n2994), .CI(\mult_827/n5 ), .CO(
        \mult_827/n4 ), .S(N6429) );
  ADDFXL \mult_827/U4  ( .A(N6419), .B(N6418), .CI(\mult_827/n4 ), .CO(
        \mult_827/n3 ), .S(N6430) );
  ADDFXL \mult_827/U3  ( .A(N6420), .B(N6419), .CI(\mult_827/n3 ), .CO(
        \mult_827/n2 ), .S(N6431) );
  ADDHXL \mult_825/U6  ( .A(N6401), .B(N6391), .CO(\mult_825/n5 ), .S(N6402)
         );
  ADDFXL \mult_825/U5  ( .A(N6392), .B(N6391), .CI(\mult_825/n5 ), .CO(
        \mult_825/n4 ), .S(N6403) );
  ADDFXL \mult_825/U4  ( .A(n2993), .B(N6392), .CI(\mult_825/n4 ), .CO(
        \mult_825/n3 ), .S(N6404) );
  ADDFXL \mult_825/U3  ( .A(N6394), .B(n2993), .CI(\mult_825/n3 ), .CO(
        \mult_825/n2 ), .S(N6405) );
  ADDHXL \mult_869/U9  ( .A(\gt_332/n9 ), .B(n3305), .CO(\mult_869/n10 ), .S(
        \mult_869/n11 ) );
  ADDHXL \mult_869/U8  ( .A(\gt_332/n15 ), .B(n3305), .CO(\mult_869/n8 ), .S(
        \mult_869/n9 ) );
  ADDHXL \mult_869/U7  ( .A(\gt_332/n9 ), .B(\gt_332/n15 ), .CO(\mult_869/n6 ), 
        .S(\mult_869/n7 ) );
  ADDHXL \mult_869/U6  ( .A(n3015), .B(\gt_332/n15 ), .CO(\mult_869/n5 ), .S(
        N6504) );
  ADDFXL \mult_869/U5  ( .A(\mult_869/n5 ), .B(n3015), .CI(\mult_869/n11 ), 
        .CO(\mult_869/n4 ), .S(N6505) );
  ADDFXL \mult_869/U4  ( .A(\mult_869/n9 ), .B(\mult_869/n10 ), .CI(
        \mult_869/n4 ), .CO(\mult_869/n3 ), .S(N6506) );
  ADDFXL \mult_869/U3  ( .A(\mult_869/n7 ), .B(\mult_869/n8 ), .CI(
        \mult_869/n3 ), .CO(\mult_869/n2 ), .S(N6507) );
  ADDFXL \mult_869/U2  ( .A(\mult_869/n6 ), .B(\gt_332/n9 ), .CI(\mult_869/n2 ), .CO(N6509), .S(N6508) );
  ADDHXL \mult_765/U6  ( .A(N5910), .B(N5926), .CO(\mult_765/n5 ), .S(N5884)
         );
  ADDFXL \mult_765/U5  ( .A(hour[2]), .B(N5926), .CI(\mult_765/n5 ), .CO(
        \mult_765/n4 ), .S(N5885) );
  ADDFXL \mult_765/U4  ( .A(hour[3]), .B(hour[2]), .CI(\mult_765/n4 ), .CO(
        \mult_765/n3 ), .S(N5886) );
  ADDFXL \mult_765/U3  ( .A(hour[4]), .B(hour[3]), .CI(\mult_765/n3 ), .CO(
        \mult_765/n2 ), .S(N5887) );
  ADDHXL \mult_769/U6  ( .A(N5910), .B(N5926), .CO(\mult_769/n5 ), .S(N5937)
         );
  ADDFXL \mult_769/U5  ( .A(n4863), .B(N5926), .CI(\mult_769/n5 ), .CO(
        \mult_769/n4 ), .S(N5938) );
  ADDFXL \mult_769/U4  ( .A(N5928), .B(n4863), .CI(\mult_769/n4 ), .CO(
        \mult_769/n3 ), .S(N5939) );
  ADDFXL \mult_769/U3  ( .A(N5929), .B(N5928), .CI(\mult_769/n3 ), .CO(
        \mult_769/n2 ), .S(N5940) );
  ADDHXL \mult_767/U6  ( .A(N5910), .B(n4858), .CO(\mult_767/n5 ), .S(N5911)
         );
  ADDFXL \mult_767/U5  ( .A(N5901), .B(n4858), .CI(\mult_767/n5 ), .CO(
        \mult_767/n4 ), .S(N5912) );
  ADDFXL \mult_767/U4  ( .A(N5902), .B(N5901), .CI(\mult_767/n4 ), .CO(
        \mult_767/n3 ), .S(N5913) );
  ADDFXL \mult_767/U3  ( .A(N5903), .B(N5902), .CI(\mult_767/n3 ), .CO(
        \mult_767/n2 ), .S(N5914) );
  ADDHXL \mult_789/U6  ( .A(N6160), .B(N6150), .CO(\mult_789/n5 ), .S(N6053)
         );
  ADDFXL \mult_789/U5  ( .A(N6151), .B(N6150), .CI(\mult_789/n5 ), .CO(
        \mult_789/n4 ), .S(N6054) );
  ADDFXL \mult_789/U4  ( .A(min[3]), .B(N6151), .CI(\mult_789/n4 ), .CO(
        \mult_789/n3 ), .S(N6055) );
  ADDFXL \mult_789/U3  ( .A(min[4]), .B(min[3]), .CI(\mult_789/n3 ), .CO(
        \mult_789/n2 ), .S(N6056) );
  ADDHXL \mult_791/U6  ( .A(N6160), .B(n4869), .CO(\mult_791/n5 ), .S(N6080)
         );
  ADDFXL \mult_791/U5  ( .A(N6070), .B(n4869), .CI(\mult_791/n5 ), .CO(
        \mult_791/n4 ), .S(N6081) );
  ADDFXL \mult_791/U4  ( .A(N6071), .B(N6070), .CI(\mult_791/n4 ), .CO(
        \mult_791/n3 ), .S(N6082) );
  ADDFXL \mult_791/U3  ( .A(N6072), .B(N6071), .CI(\mult_791/n3 ), .CO(
        \mult_791/n2 ), .S(N6083) );
  ADDHXL \mult_793/U6  ( .A(N6160), .B(N6150), .CO(\mult_793/n5 ), .S(N6107)
         );
  ADDFXL \mult_793/U5  ( .A(n4867), .B(N6150), .CI(\mult_793/n5 ), .CO(
        \mult_793/n4 ), .S(N6108) );
  ADDFXL \mult_793/U4  ( .A(N6098), .B(n4867), .CI(\mult_793/n4 ), .CO(
        \mult_793/n3 ), .S(N6109) );
  ADDFXL \mult_793/U3  ( .A(N6099), .B(N6098), .CI(\mult_793/n3 ), .CO(
        \mult_793/n2 ), .S(N6110) );
  ADDHXL \mult_795/U6  ( .A(N6160), .B(n4869), .CO(\mult_795/n5 ), .S(N6134)
         );
  ADDFXL \mult_795/U5  ( .A(N6124), .B(n4869), .CI(\mult_795/n5 ), .CO(
        \mult_795/n4 ), .S(N6135) );
  ADDFXL \mult_795/U4  ( .A(N6125), .B(N6124), .CI(\mult_795/n4 ), .CO(
        \mult_795/n3 ), .S(N6136) );
  ADDFXL \mult_795/U3  ( .A(N6126), .B(N6125), .CI(\mult_795/n3 ), .CO(
        \mult_795/n2 ), .S(N6137) );
  ADDHXL \mult_799/U6  ( .A(N6160), .B(n4869), .CO(\mult_799/n5 ), .S(N6187)
         );
  ADDFXL \mult_799/U5  ( .A(N6177), .B(n4869), .CI(\mult_799/n5 ), .CO(
        \mult_799/n4 ), .S(N6188) );
  ADDFXL \mult_799/U4  ( .A(N6178), .B(N6177), .CI(\mult_799/n4 ), .CO(
        \mult_799/n3 ), .S(N6189) );
  ADDFXL \mult_799/U3  ( .A(N6179), .B(N6178), .CI(\mult_799/n3 ), .CO(
        \mult_799/n2 ), .S(N6190) );
  ADDHXL \mult_797/U6  ( .A(N6160), .B(N6150), .CO(\mult_797/n5 ), .S(N6161)
         );
  ADDFXL \mult_797/U5  ( .A(N6151), .B(N6150), .CI(\mult_797/n5 ), .CO(
        \mult_797/n4 ), .S(N6162) );
  ADDFXL \mult_797/U4  ( .A(n4868), .B(N6151), .CI(\mult_797/n4 ), .CO(
        \mult_797/n3 ), .S(N6163) );
  ADDFXL \mult_797/U3  ( .A(N6153), .B(n4868), .CI(\mult_797/n3 ), .CO(
        \mult_797/n2 ), .S(N6164) );
  DFFRX1 \cycle_reg[0]  ( .D(cycle_n[0]), .CK(clk), .RN(n3127), .Q(cycle[0]), 
        .QN(n4744) );
  DFFRX1 \cycle_reg[9]  ( .D(cycle_n[9]), .CK(clk), .RN(n3124), .Q(cycle[9]), 
        .QN(n4694) );
  DFFRX1 \cycle_reg[1]  ( .D(cycle_n[1]), .CK(clk), .RN(n3124), .Q(cycle[1]), 
        .QN(n4745) );
  DFFRX1 \cycle_reg[2]  ( .D(cycle_n[2]), .CK(clk), .RN(n3124), .Q(cycle[2]), 
        .QN(n4689) );
  DFFRX1 \cycle_reg[3]  ( .D(cycle_n[3]), .CK(clk), .RN(n3124), .Q(cycle[3]), 
        .QN(n4690) );
  DFFRX1 \cycle_reg[4]  ( .D(cycle_n[4]), .CK(clk), .RN(n3124), .Q(cycle[4]), 
        .QN(n4691) );
  DFFRX1 \cycle_reg[5]  ( .D(cycle_n[5]), .CK(clk), .RN(n3124), .Q(cycle[5]), 
        .QN(n4692) );
  DFFRX1 \cycle_reg[6]  ( .D(cycle_n[6]), .CK(clk), .RN(n3124), .Q(cycle[6]), 
        .QN(n4701) );
  DFFRX1 \cycle_reg[7]  ( .D(cycle_n[7]), .CK(clk), .RN(n3124), .Q(cycle[7]), 
        .QN(n4693) );
  DFFRX1 \cycle_reg[8]  ( .D(cycle_n[8]), .CK(clk), .RN(n3124), .Q(cycle[8]), 
        .QN(n4702) );
  DFFRX1 \cycle_reg[10]  ( .D(cycle_n[10]), .CK(clk), .RN(n3125), .Q(cycle[10]), .QN(n4703) );
  DFFRX1 \cycle_reg[11]  ( .D(cycle_n[11]), .CK(clk), .RN(n3125), .Q(cycle[11]), .QN(n4704) );
  DFFRX1 \cycle_reg[12]  ( .D(cycle_n[12]), .CK(clk), .RN(n3125), .Q(cycle[12]), .QN(n4695) );
  DFFRX1 \cycle_reg[13]  ( .D(cycle_n[13]), .CK(clk), .RN(n3125), .Q(cycle[13]), .QN(n4696) );
  DFFRX1 \cycle_reg[14]  ( .D(cycle_n[14]), .CK(clk), .RN(n3125), .Q(cycle[14]), .QN(n4697) );
  DFFRX1 \cycle_reg[15]  ( .D(cycle_n[15]), .CK(clk), .RN(n3125), .Q(cycle[15]), .QN(n4698) );
  DFFRX1 \cycle_reg[16]  ( .D(cycle_n[16]), .CK(clk), .RN(n3125), .Q(cycle[16]), .QN(n4705) );
  DFFRX1 \cycle_reg[17]  ( .D(cycle_n[17]), .CK(clk), .RN(n3124), .Q(cycle[17]), .QN(n4706) );
  DFFRX1 \cycle_reg[18]  ( .D(cycle_n[18]), .CK(clk), .RN(n3124), .Q(cycle[18]), .QN(n4700) );
  DFFRX1 \cycle_reg[19]  ( .D(cycle_n[19]), .CK(clk), .RN(n3124), .Q(cycle[19]), .QN(n4699) );
  DFFRX2 \hour_reg[1]  ( .D(hour_n[1]), .CK(clk), .RN(n3125), .Q(N5926), .QN(
        n4858) );
  DFFRX2 \hour_reg[3]  ( .D(hour_n[3]), .CK(clk), .RN(n3134), .Q(hour[3]), 
        .QN(n4862) );
  DFFRX1 \hour_reg[5]  ( .D(hour_n[5]), .CK(clk), .RN(n3124), .Q(hour[5]), 
        .QN(n4859) );
  DFFRX1 \hour_reg[6]  ( .D(hour_n[6]), .CK(clk), .RN(n3133), .Q(hour[6]), 
        .QN(n4860) );
  DFFRX1 \min_reg[6]  ( .D(min_n[6]), .CK(clk), .RN(n3126), .Q(min[6]), .QN(
        n4865) );
  XOR3XL \add_769/U1_8  ( .A(N5941), .B(n3073), .C(\add_769/carry[8] ), .Y(
        N5950) );
  XOR3XL \add_767/U1_8  ( .A(N5915), .B(n3073), .C(\add_767/carry[8] ), .Y(
        N5924) );
  XOR3XL \add_765/U1_8  ( .A(N5888), .B(n3073), .C(\add_765/carry[8] ), .Y(
        N5897) );
  XOR3XL \add_799/U1_8  ( .A(N6191), .B(n3073), .C(\add_799/carry[8] ), .Y(
        N6200) );
  XOR3XL \add_827/U1_8  ( .A(N6432), .B(n3073), .C(\add_827/carry[8] ), .Y(
        N6441) );
  XOR3XL \add_0_root_add_0_root_add_609_4_cf/U1_19  ( .A(N7686), .B(N4433), 
        .C(\add_0_root_add_0_root_add_609_4_cf/carry[19] ), .Y(N4473) );
  XOR3XL \add_0_root_add_0_root_add_579_4_cf/U1_19  ( .A(N7666), .B(N668), .C(
        \add_0_root_add_0_root_add_579_4_cf/carry[19] ), .Y(N4195) );
  XOR3XL \add_0_root_add_0_root_add_601_3/U1_19  ( .A(N4343), .B(N4323), .C(
        \add_0_root_add_0_root_add_601_3/carry[19] ), .Y(N4383) );
  XOR3XL \add_0_root_add_0_root_add_661_4_cf/U1_19  ( .A(N7604), .B(N668), .C(
        \add_0_root_add_0_root_add_661_4_cf/carry[19] ), .Y(N5040) );
  ADDFXL \add_765/U1_4  ( .A(N5884), .B(n3075), .CI(n2960), .CO(
        \add_765/carry[5] ), .S(N5893) );
  ADDFXL \add_767/U1_4  ( .A(N5911), .B(n3075), .CI(n2960), .CO(
        \add_767/carry[5] ), .S(N5920) );
  ADDFXL \add_769/U1_4  ( .A(N5937), .B(n3075), .CI(n2960), .CO(
        \add_769/carry[5] ), .S(N5946) );
  ADDFXL \add_799/U1_4  ( .A(N6187), .B(n3075), .CI(n2954), .CO(
        \add_799/carry[5] ), .S(N6196) );
  ADDFXL \add_797/U1_4  ( .A(N6161), .B(n3075), .CI(n2954), .CO(
        \add_797/carry[5] ), .S(N6170) );
  ADDFXL \add_795/U1_4  ( .A(N6134), .B(n3075), .CI(n2954), .CO(
        \add_795/carry[5] ), .S(N6143) );
  ADDFXL \add_789/U1_4  ( .A(N6053), .B(n3075), .CI(n2954), .CO(
        \add_789/carry[5] ), .S(N6062) );
  ADDFXL \add_791/U1_4  ( .A(N6080), .B(n3075), .CI(n2954), .CO(
        \add_791/carry[5] ), .S(N6089) );
  ADDFXL \add_793/U1_4  ( .A(N6107), .B(n3075), .CI(n2954), .CO(
        \add_793/carry[5] ), .S(N6116) );
  ADDFXL \add_827/U1_4  ( .A(N6428), .B(n3075), .CI(n2955), .CO(
        \add_827/carry[5] ), .S(N6437) );
  ADDFXL \add_825/U1_4  ( .A(N6402), .B(n3075), .CI(n2955), .CO(
        \add_825/carry[5] ), .S(N6411) );
  ADDFXL \add_823/U1_4  ( .A(N6375), .B(n3075), .CI(n2955), .CO(
        \add_823/carry[5] ), .S(N6384) );
  ADDFXL \add_817/U1_4  ( .A(N6294), .B(n3075), .CI(n2955), .CO(
        \add_817/carry[5] ), .S(N6303) );
  ADDFXL \add_819/U1_4  ( .A(N6321), .B(n3075), .CI(n2955), .CO(
        \add_819/carry[5] ), .S(N6330) );
  ADDFXL \add_821/U1_4  ( .A(N6348), .B(n3075), .CI(n2955), .CO(
        \add_821/carry[5] ), .S(N6357) );
  ADDFXL \add_765/U1_5  ( .A(N5885), .B(n3081), .CI(\add_765/carry[5] ), .CO(
        \add_765/carry[6] ), .S(N5894) );
  ADDFXL \add_767/U1_5  ( .A(N5912), .B(n3081), .CI(\add_767/carry[5] ), .CO(
        \add_767/carry[6] ), .S(N5921) );
  ADDFXL \add_769/U1_5  ( .A(N5938), .B(n3081), .CI(\add_769/carry[5] ), .CO(
        \add_769/carry[6] ), .S(N5947) );
  ADDFXL \add_765/U1_6  ( .A(N5886), .B(n3077), .CI(\add_765/carry[6] ), .CO(
        \add_765/carry[7] ), .S(N5895) );
  ADDFXL \add_767/U1_6  ( .A(N5913), .B(n3077), .CI(\add_767/carry[6] ), .CO(
        \add_767/carry[7] ), .S(N5922) );
  ADDFXL \add_769/U1_6  ( .A(N5939), .B(n3077), .CI(\add_769/carry[6] ), .CO(
        \add_769/carry[7] ), .S(N5948) );
  ADDFXL \add_799/U1_6  ( .A(N6189), .B(n3077), .CI(\add_799/carry[6] ), .CO(
        \add_799/carry[7] ), .S(N6198) );
  ADDFXL \add_797/U1_6  ( .A(N6163), .B(n3077), .CI(\add_797/carry[6] ), .CO(
        \add_797/carry[7] ), .S(N6172) );
  ADDFXL \add_795/U1_6  ( .A(N6136), .B(n3077), .CI(\add_795/carry[6] ), .CO(
        \add_795/carry[7] ), .S(N6145) );
  ADDFXL \add_789/U1_6  ( .A(N6055), .B(n3077), .CI(\add_789/carry[6] ), .CO(
        \add_789/carry[7] ), .S(N6064) );
  ADDFXL \add_791/U1_6  ( .A(N6082), .B(n3077), .CI(\add_791/carry[6] ), .CO(
        \add_791/carry[7] ), .S(N6091) );
  ADDFXL \add_793/U1_6  ( .A(N6109), .B(n3077), .CI(\add_793/carry[6] ), .CO(
        \add_793/carry[7] ), .S(N6118) );
  ADDFXL \add_827/U1_6  ( .A(N6430), .B(n3077), .CI(\add_827/carry[6] ), .CO(
        \add_827/carry[7] ), .S(N6439) );
  ADDFXL \add_825/U1_6  ( .A(N6404), .B(n3077), .CI(\add_825/carry[6] ), .CO(
        \add_825/carry[7] ), .S(N6413) );
  ADDFXL \add_823/U1_6  ( .A(N6377), .B(n3077), .CI(\add_823/carry[6] ), .CO(
        \add_823/carry[7] ), .S(N6386) );
  ADDFXL \add_817/U1_6  ( .A(N6296), .B(n3077), .CI(\add_817/carry[6] ), .CO(
        \add_817/carry[7] ), .S(N6305) );
  ADDFXL \add_819/U1_6  ( .A(N6323), .B(n3077), .CI(\add_819/carry[6] ), .CO(
        \add_819/carry[7] ), .S(N6332) );
  ADDFXL \add_821/U1_6  ( .A(N6350), .B(n3077), .CI(\add_821/carry[6] ), .CO(
        \add_821/carry[7] ), .S(N6359) );
  ADDFXL \add_765/U1_7  ( .A(N5887), .B(n3079), .CI(\add_765/carry[7] ), .CO(
        \add_765/carry[8] ), .S(N5896) );
  ADDFXL \add_767/U1_7  ( .A(N5914), .B(n3079), .CI(\add_767/carry[7] ), .CO(
        \add_767/carry[8] ), .S(N5923) );
  ADDFXL \add_769/U1_7  ( .A(N5940), .B(n3079), .CI(\add_769/carry[7] ), .CO(
        \add_769/carry[8] ), .S(N5949) );
  ADDFXL \add_799/U1_7  ( .A(N6190), .B(n3079), .CI(\add_799/carry[7] ), .CO(
        \add_799/carry[8] ), .S(N6199) );
  ADDFXL \add_797/U1_7  ( .A(N6164), .B(n3079), .CI(\add_797/carry[7] ), .CO(
        \add_797/carry[8] ), .S(N6173) );
  ADDFXL \add_795/U1_7  ( .A(N6137), .B(n3079), .CI(\add_795/carry[7] ), .CO(
        \add_795/carry[8] ), .S(N6146) );
  ADDFXL \add_789/U1_7  ( .A(N6056), .B(n3079), .CI(\add_789/carry[7] ), .CO(
        \add_789/carry[8] ), .S(N6065) );
  ADDFXL \add_791/U1_7  ( .A(N6083), .B(n3079), .CI(\add_791/carry[7] ), .CO(
        \add_791/carry[8] ), .S(N6092) );
  ADDFXL \add_793/U1_7  ( .A(N6110), .B(n3079), .CI(\add_793/carry[7] ), .CO(
        \add_793/carry[8] ), .S(N6119) );
  ADDFXL \add_827/U1_7  ( .A(N6431), .B(n3079), .CI(\add_827/carry[7] ), .CO(
        \add_827/carry[8] ), .S(N6440) );
  ADDFXL \add_825/U1_7  ( .A(N6405), .B(n3079), .CI(\add_825/carry[7] ), .CO(
        \add_825/carry[8] ), .S(N6414) );
  ADDFXL \add_823/U1_7  ( .A(N6378), .B(n3079), .CI(\add_823/carry[7] ), .CO(
        \add_823/carry[8] ), .S(N6387) );
  ADDFXL \add_817/U1_7  ( .A(N6297), .B(n3079), .CI(\add_817/carry[7] ), .CO(
        \add_817/carry[8] ), .S(N6306) );
  ADDFXL \add_819/U1_7  ( .A(N6324), .B(n3079), .CI(\add_819/carry[7] ), .CO(
        \add_819/carry[8] ), .S(N6333) );
  ADDFXL \add_821/U1_7  ( .A(N6351), .B(n3079), .CI(\add_821/carry[7] ), .CO(
        \add_821/carry[8] ), .S(N6360) );
  XOR3XL \add_797/U1_8  ( .A(N6165), .B(n3073), .C(\add_797/carry[8] ), .Y(
        N6174) );
  XOR3XL \add_795/U1_8  ( .A(N6138), .B(n3073), .C(\add_795/carry[8] ), .Y(
        N6147) );
  XOR3XL \add_789/U1_8  ( .A(N6057), .B(n3073), .C(\add_789/carry[8] ), .Y(
        N6066) );
  XOR3XL \add_791/U1_8  ( .A(N6084), .B(n3073), .C(\add_791/carry[8] ), .Y(
        N6093) );
  XOR3XL \add_793/U1_8  ( .A(N6111), .B(n3073), .C(\add_793/carry[8] ), .Y(
        N6120) );
  XOR3XL \add_825/U1_8  ( .A(N6406), .B(n3073), .C(\add_825/carry[8] ), .Y(
        N6415) );
  XOR3XL \add_823/U1_8  ( .A(N6379), .B(n3073), .C(\add_823/carry[8] ), .Y(
        N6388) );
  XOR3XL \add_817/U1_8  ( .A(N6298), .B(n3073), .C(\add_817/carry[8] ), .Y(
        N6307) );
  XOR3XL \add_819/U1_8  ( .A(N6325), .B(n3073), .C(\add_819/carry[8] ), .Y(
        N6334) );
  XOR3XL \add_821/U1_8  ( .A(N6352), .B(n3073), .C(\add_821/carry[8] ), .Y(
        N6361) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_3  ( .A(N7702), .B(N4431), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[3] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[4] ), .S(N4457) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_3  ( .A(N4327), .B(n4856), .CI(
        \add_0_root_add_0_root_add_601_3/carry[3] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[4] ), .S(N4367) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_4  ( .A(N673), .B(N667), .CI(
        \add_0_root_add_0_root_add_209_3/carry[4] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[5] ), .S(N713) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_4  ( .A(N1385), .B(N667), .CI(
        \add_0_root_add_1_root_add_282_4/carry[4] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[5] ), .S(N1445) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_4  ( .A(N7701), .B(N4432), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[4] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[5] ), .S(N4458) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_4  ( .A(N7681), .B(N667), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[4] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[5] ), .S(N4180) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_4  ( .A(N4328), .B(N4322), .CI(
        \add_0_root_add_0_root_add_601_3/carry[4] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[5] ), .S(N4368) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_5  ( .A(N674), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[5] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[6] ), .S(N714) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_5  ( .A(N1386), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[5] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[6] ), .S(N1446) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_6  ( .A(N675), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[6] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[7] ), .S(N715) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_6  ( .A(N1387), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[6] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[7] ), .S(N1447) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_7  ( .A(N676), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[7] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[8] ), .S(N716) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_7  ( .A(N1388), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[7] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[8] ), .S(N1448) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_8  ( .A(N7697), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[8] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[9] ), .S(N4462) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_8  ( .A(N4332), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[8] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[9] ), .S(N4372) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_8  ( .A(N7677), .B(N668), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[8] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[9] ), .S(N4184) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_8  ( .A(N677), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[8] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[9] ), .S(N717) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_8  ( .A(N1389), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[8] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[9] ), .S(N1449) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_9  ( .A(N7696), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[9] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[10] ), .S(N4463) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_9  ( .A(N4333), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[9] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[10] ), .S(N4373) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_9  ( .A(N7676), .B(N668), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[9] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[10] ), .S(N4185) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_9  ( .A(N678), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[9] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[10] ), .S(N718) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_9  ( .A(N1390), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[9] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[10] ), .S(N1450) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_10  ( .A(N7695), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[10] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[11] ), .S(N4464) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_10  ( .A(N4334), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[10] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[11] ), .S(N4374) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_10  ( .A(N7675), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[10] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[11] ), .S(N4186) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_10  ( .A(N679), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[10] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[11] ), .S(N719) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_10  ( .A(N1391), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[10] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[11] ), .S(N1451) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_11  ( .A(N7694), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[11] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[12] ), .S(N4465) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_11  ( .A(N4335), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[11] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[12] ), .S(N4375) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_11  ( .A(N7674), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[11] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[12] ), .S(N4187) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_11  ( .A(N680), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[11] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[12] ), .S(N720) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_11  ( .A(N1392), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[11] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[12] ), .S(N1452) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_12  ( .A(N7693), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[12] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[13] ), .S(N4466) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_12  ( .A(N4336), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[12] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[13] ), .S(N4376) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_12  ( .A(N7673), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[12] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[13] ), .S(N4188) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_12  ( .A(N681), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[12] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[13] ), .S(N721) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_12  ( .A(N1393), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[12] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[13] ), .S(N1453) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_13  ( .A(N7692), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[13] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[14] ), .S(N4467) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_13  ( .A(N4337), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[13] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[14] ), .S(N4377) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_13  ( .A(N7672), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[13] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[14] ), .S(N4189) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_13  ( .A(N682), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[13] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[14] ), .S(N722) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_13  ( .A(N1394), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[13] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[14] ), .S(N1454) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_14  ( .A(N7691), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[14] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[15] ), .S(N4468) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_14  ( .A(N4338), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[14] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[15] ), .S(N4378) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_14  ( .A(N7671), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[14] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[15] ), .S(N4190) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_14  ( .A(N683), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[14] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[15] ), .S(N723) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_14  ( .A(N1395), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[14] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[15] ), .S(N1455) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_15  ( .A(N7690), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[15] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[16] ), .S(N4469) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_15  ( .A(N4339), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[15] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[16] ), .S(N4379) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_15  ( .A(N7670), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[15] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[16] ), .S(N4191) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_15  ( .A(N684), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[15] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[16] ), .S(N724) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_15  ( .A(N1396), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[15] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[16] ), .S(N1456) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_16  ( .A(N7689), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[16] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[17] ), .S(N4470) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_16  ( .A(N4340), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[16] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[17] ), .S(N4380) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_16  ( .A(N7669), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[16] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[17] ), .S(N4192) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_16  ( .A(N685), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[16] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[17] ), .S(N725) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_16  ( .A(N1397), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[16] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[17] ), .S(N1457) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_17  ( .A(N7688), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[17] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[18] ), .S(N4471) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_17  ( .A(N4341), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[17] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[18] ), .S(N4381) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_17  ( .A(N7668), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[17] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[18] ), .S(N4193) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_17  ( .A(N686), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[17] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[18] ), .S(N726) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_17  ( .A(N1398), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[17] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[18] ), .S(N1458) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_18  ( .A(N7687), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[18] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[19] ), .S(N4472) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_18  ( .A(N4342), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[18] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[19] ), .S(N4382) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_18  ( .A(N7667), .B(N668), 
        .CI(\add_0_root_add_0_root_add_579_4_cf/carry[18] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[19] ), .S(N4194) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_18  ( .A(N687), .B(N668), .CI(
        \add_0_root_add_0_root_add_209_3/carry[18] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[19] ), .S(N727) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_18  ( .A(N1399), .B(N668), .CI(
        \add_0_root_add_1_root_add_282_4/carry[18] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[19] ), .S(N1459) );
  XOR3XL \add_0_root_add_0_root_add_446_3/U1_19  ( .A(N2829), .B(N668), .C(
        \add_0_root_add_0_root_add_446_3/carry[19] ), .Y(N2869) );
  XOR3XL \add_0_root_add_0_root_add_209_3/U1_19  ( .A(N688), .B(N668), .C(
        \add_0_root_add_0_root_add_209_3/carry[19] ), .Y(N728) );
  XOR3XL \add_0_root_add_1_root_add_282_4/U1_19  ( .A(N1400), .B(N668), .C(
        \add_0_root_add_1_root_add_282_4/carry[19] ), .Y(N1460) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_18  ( .A(N7605), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[18] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[19] ), .S(N5039) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_2  ( .A(N7703), .B(n4855), 
        .CI(n2962), .CO(\add_0_root_add_0_root_add_609_4_cf/carry[3] ), .S(
        N4456) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_2  ( .A(N4326), .B(n3305), .CI(
        n2971), .CO(\add_0_root_add_0_root_add_601_3/carry[3] ), .S(N4366) );
  ADDFXL \add_799/U1_5  ( .A(N6188), .B(n3081), .CI(\add_799/carry[5] ), .CO(
        \add_799/carry[6] ), .S(N6197) );
  ADDFXL \add_797/U1_5  ( .A(N6162), .B(n3081), .CI(\add_797/carry[5] ), .CO(
        \add_797/carry[6] ), .S(N6171) );
  ADDFXL \add_795/U1_5  ( .A(N6135), .B(n3081), .CI(\add_795/carry[5] ), .CO(
        \add_795/carry[6] ), .S(N6144) );
  ADDFXL \add_789/U1_5  ( .A(N6054), .B(n3081), .CI(\add_789/carry[5] ), .CO(
        \add_789/carry[6] ), .S(N6063) );
  ADDFXL \add_791/U1_5  ( .A(N6081), .B(n3081), .CI(\add_791/carry[5] ), .CO(
        \add_791/carry[6] ), .S(N6090) );
  ADDFXL \add_793/U1_5  ( .A(N6108), .B(n3081), .CI(\add_793/carry[5] ), .CO(
        \add_793/carry[6] ), .S(N6117) );
  ADDFXL \add_827/U1_5  ( .A(N6429), .B(n3081), .CI(\add_827/carry[5] ), .CO(
        \add_827/carry[6] ), .S(N6438) );
  ADDFXL \add_825/U1_5  ( .A(N6403), .B(n3081), .CI(\add_825/carry[5] ), .CO(
        \add_825/carry[6] ), .S(N6412) );
  ADDFXL \add_823/U1_5  ( .A(N6376), .B(n3081), .CI(\add_823/carry[5] ), .CO(
        \add_823/carry[6] ), .S(N6385) );
  ADDFXL \add_817/U1_5  ( .A(N6295), .B(n3081), .CI(\add_817/carry[5] ), .CO(
        \add_817/carry[6] ), .S(N6304) );
  ADDFXL \add_819/U1_5  ( .A(N6322), .B(n3081), .CI(\add_819/carry[5] ), .CO(
        \add_819/carry[6] ), .S(N6331) );
  ADDFXL \add_821/U1_5  ( .A(N6349), .B(n3081), .CI(\add_821/carry[5] ), .CO(
        \add_821/carry[6] ), .S(N6358) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_3  ( .A(N7620), .B(N666), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[3] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[4] ), .S(N5024) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_4  ( .A(N2814), .B(N667), .CI(
        \add_0_root_add_0_root_add_446_3/carry[4] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[5] ), .S(N2854) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_4  ( .A(N7619), .B(N667), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[4] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[5] ), .S(N5025) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_5  ( .A(N4329), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[5] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[6] ), .S(N4369) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_5  ( .A(N7700), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[5] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[6] ), .S(N4459) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_5  ( .A(N7680), .B(N668), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[5] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[6] ), .S(N4181) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_5  ( .A(N2815), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[5] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[6] ), .S(N2855) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_6  ( .A(N4330), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[6] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[7] ), .S(N4370) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_6  ( .A(N7699), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[6] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[7] ), .S(N4460) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_6  ( .A(N7679), .B(N668), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[6] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[7] ), .S(N4182) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_6  ( .A(N2816), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[6] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[7] ), .S(N2856) );
  ADDFXL \add_0_root_add_0_root_add_601_3/U1_7  ( .A(N4331), .B(N4323), .CI(
        \add_0_root_add_0_root_add_601_3/carry[7] ), .CO(
        \add_0_root_add_0_root_add_601_3/carry[8] ), .S(N4371) );
  ADDFXL \add_0_root_add_0_root_add_609_4_cf/U1_7  ( .A(N7698), .B(N4433), 
        .CI(\add_0_root_add_0_root_add_609_4_cf/carry[7] ), .CO(
        \add_0_root_add_0_root_add_609_4_cf/carry[8] ), .S(N4461) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_7  ( .A(N7678), .B(N668), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[7] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[8] ), .S(N4183) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_7  ( .A(N2817), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[7] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[8] ), .S(N2857) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_8  ( .A(N2818), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[8] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[9] ), .S(N2858) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_8  ( .A(N7615), .B(N668), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[8] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[9] ), .S(N5029) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_9  ( .A(N2819), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[9] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[10] ), .S(N2859) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_9  ( .A(N7614), .B(N668), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[9] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[10] ), .S(N5030) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_10  ( .A(N2820), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[10] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[11] ), .S(N2860) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_10  ( .A(N7613), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[10] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[11] ), .S(N5031) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_11  ( .A(N2821), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[11] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[12] ), .S(N2861) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_12  ( .A(N2822), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[12] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[13] ), .S(N2862) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_12  ( .A(N7611), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[12] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[13] ), .S(N5033) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_13  ( .A(N2823), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[13] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[14] ), .S(N2863) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_13  ( .A(N7610), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[13] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[14] ), .S(N5034) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_14  ( .A(N2824), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[14] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[15] ), .S(N2864) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_15  ( .A(N2825), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[15] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[16] ), .S(N2865) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_16  ( .A(N2826), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[16] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[17] ), .S(N2866) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_17  ( .A(N2827), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[17] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[18] ), .S(N2867) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_17  ( .A(N7606), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[17] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[18] ), .S(N5038) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_18  ( .A(N2828), .B(N668), .CI(
        \add_0_root_add_0_root_add_446_3/carry[18] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[19] ), .S(N2868) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_2  ( .A(N7621), .B(n4855), 
        .CI(n2970), .CO(\add_0_root_add_0_root_add_661_4_cf/carry[3] ), .S(
        N5023) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_2  ( .A(N2812), .B(n4855), .CI(
        n2969), .CO(\add_0_root_add_0_root_add_446_3/carry[3] ), .S(N2852) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_5  ( .A(N7618), .B(N668), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[5] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[6] ), .S(N5026) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_6  ( .A(N7617), .B(N668), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[6] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[7] ), .S(N5027) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_7  ( .A(N7616), .B(N668), .CI(
        \add_0_root_add_0_root_add_661_4_cf/carry[7] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[8] ), .S(N5028) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_11  ( .A(N7612), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[11] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[12] ), .S(N5032) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_14  ( .A(N7609), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[14] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[15] ), .S(N5035) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_15  ( .A(N7608), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[15] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[16] ), .S(N5036) );
  ADDFXL \add_0_root_add_0_root_add_661_4_cf/U1_16  ( .A(N7607), .B(N668), 
        .CI(\add_0_root_add_0_root_add_661_4_cf/carry[16] ), .CO(
        \add_0_root_add_0_root_add_661_4_cf/carry[17] ), .S(N5037) );
  DFFRX4 \offset_reg[9]  ( .D(n1646), .CK(clk), .RN(n3134), .Q(N798), .QN(
        n2986) );
  DFFRX4 \FB_A_reg[18]  ( .D(n1612), .CK(clk), .RN(n3129), .Q(N4427), .QN(
        n4799) );
  DFFRX4 \sec_reg[1]  ( .D(n1620), .CK(clk), .RN(n3141), .Q(N6391), .QN(n2994)
         );
  DFFRX4 \FB_A_reg[2]  ( .D(n1596), .CK(clk), .RN(n3130), .Q(N4411), .QN(n4796) );
  DFFRX2 \pix_c_reg[3]  ( .D(n1664), .CK(clk), .RN(n3127), .Q(\gt_332/n9 ), 
        .QN(n4857) );
  DFFRX2 \offset_w_reg[7]  ( .D(n1631), .CK(clk), .RN(n3138), .Q(N4352), .QN(
        n4730) );
  DFFRX2 \pic_A_reg[0]  ( .D(n1444), .CK(clk), .RN(n3124), .Q(pic_A[0]), .QN(
        n4727) );
  DFFRX4 \pix_c_reg[2]  ( .D(n1679), .CK(clk), .RN(n3127), .Q(\gt_332/n15 ), 
        .QN(n4856) );
  DFFRX4 \sec_reg[3]  ( .D(n1622), .CK(clk), .RN(n3141), .Q(sec[3]), .QN(n2993) );
  DFFRX2 \pic_A_reg[5]  ( .D(n1449), .CK(clk), .RN(n3136), .Q(pic_A[5]), .QN(
        n4712) );
  DFFRX4 \FB_A_reg[0]  ( .D(n1594), .CK(clk), .RN(n3130), .Q(N4409), .QN(n4808) );
  DFFRX2 \pic_A_reg[1]  ( .D(n1445), .CK(clk), .RN(n3133), .Q(pic_A[1]), .QN(
        n4716) );
  DFFRX4 \offset_reg[10]  ( .D(n1652), .CK(clk), .RN(n3138), .Q(N799), .QN(
        n2987) );
  DFFRX4 \FB_A_reg[17]  ( .D(n1611), .CK(clk), .RN(n3129), .Q(N4426), .QN(
        n4800) );
  DFFRX4 \FB_A_reg[8]  ( .D(n1602), .CK(clk), .RN(n3130), .Q(N4417), .QN(n4790) );
  DFFRX4 \FB_A_reg[16]  ( .D(n1610), .CK(clk), .RN(n3129), .Q(N4425), .QN(
        n4801) );
  DFFRX4 \FB_A_reg[10]  ( .D(n1604), .CK(clk), .RN(n3130), .Q(N4419), .QN(
        n4807) );
  DFFRX4 \FB_A_reg[11]  ( .D(n1605), .CK(clk), .RN(n3130), .Q(N4420), .QN(
        n4806) );
  DFFRX4 \FB_A_reg[13]  ( .D(n1607), .CK(clk), .RN(n3129), .Q(N4422), .QN(
        n4804) );
  DFFRX4 \FB_A_reg[14]  ( .D(n1608), .CK(clk), .RN(n3129), .Q(N4423), .QN(
        n4803) );
  DFFRX4 \FB_A_reg[15]  ( .D(n1609), .CK(clk), .RN(n3129), .Q(N4424), .QN(
        n4802) );
  DFFRX4 \sec_reg[2]  ( .D(n1621), .CK(clk), .RN(n3141), .Q(N6392), .QN(n2995)
         );
  DFFRX4 \offset_w_reg[0]  ( .D(n1677), .CK(clk), .RN(n3137), .Q(N4345), .QN(
        n4743) );
  DFFRX4 \FB_A_reg[5]  ( .D(n1599), .CK(clk), .RN(n3130), .Q(N4414), .QN(n4793) );
  DFFRX4 \FB_A_reg[6]  ( .D(n1600), .CK(clk), .RN(n3138), .Q(N4415), .QN(n4792) );
  DFFRX4 \FB_A_reg[7]  ( .D(n1601), .CK(clk), .RN(n3130), .Q(N4416), .QN(n4791) );
  DFFRX4 \FB_A_reg[3]  ( .D(n1597), .CK(clk), .RN(n3130), .Q(N4412), .QN(n4795) );
  DFFRX4 \FB_A_reg[4]  ( .D(n1598), .CK(clk), .RN(n3130), .Q(N4413), .QN(n4794) );
  DFFRX2 \FB_A_reg[19]  ( .D(n1613), .CK(clk), .RN(n3129), .Q(N4428), .QN(
        n4798) );
  DFFRX2 \pic_A_reg[18]  ( .D(n1462), .CK(clk), .RN(n3131), .Q(pic_A[18]), 
        .QN(n4718) );
  DFFRX2 \pic_A_reg[16]  ( .D(n1460), .CK(clk), .RN(n3131), .Q(pic_A[16]), 
        .QN(n4720) );
  DFFRX2 \pic_A_reg[17]  ( .D(n1461), .CK(clk), .RN(n3131), .Q(pic_A[17]), 
        .QN(n4719) );
  DFFRX2 \pic_A_reg[6]  ( .D(n1450), .CK(clk), .RN(n3126), .Q(pic_A[6]), .QN(
        n4711) );
  DFFRX2 \pic_A_reg[7]  ( .D(n1451), .CK(clk), .RN(n3124), .Q(pic_A[7]), .QN(
        n4710) );
  DFFRX2 \pic_A_reg[8]  ( .D(n1452), .CK(clk), .RN(n3136), .Q(pic_A[8]), .QN(
        n4709) );
  DFFRX2 \pic_A_reg[9]  ( .D(n1453), .CK(clk), .RN(n3124), .Q(pic_A[9]), .QN(
        n4708) );
  DFFRX2 \pic_A_reg[11]  ( .D(n1455), .CK(clk), .RN(n3140), .Q(pic_A[11]), 
        .QN(n4725) );
  DFFRX2 \pic_A_reg[13]  ( .D(n1457), .CK(clk), .RN(n3124), .Q(pic_A[13]), 
        .QN(n4723) );
  DFFRX2 \pic_A_reg[14]  ( .D(n1458), .CK(clk), .RN(n3131), .Q(pic_A[14]), 
        .QN(n4722) );
  DFFRX2 \pic_A_reg[15]  ( .D(n1459), .CK(clk), .RN(n3131), .Q(pic_A[15]), 
        .QN(n4721) );
  DFFRX2 \sec_reg[5]  ( .D(n1624), .CK(clk), .RN(n3135), .Q(sec[5]), .QN(n3115) );
  DFFRX4 \offset_reg[11]  ( .D(n1647), .CK(clk), .RN(n3141), .Q(N800), .QN(
        n2988) );
  DFFRX4 \FB_A_reg[12]  ( .D(n1606), .CK(clk), .RN(n3129), .Q(N4421), .QN(
        n4805) );
  DFFRX4 \FB_A_reg[9]  ( .D(n1603), .CK(clk), .RN(n3130), .Q(N4418), .QN(n4789) );
  DFFRX4 \sec_reg[4]  ( .D(n1623), .CK(clk), .RN(n3136), .Q(sec[4]), .QN(n2977) );
  DFFRX2 \pic_A_reg[10]  ( .D(n1454), .CK(clk), .RN(n3136), .Q(pic_A[10]), 
        .QN(n4726) );
  DFFRX2 \pic_A_reg[12]  ( .D(n1456), .CK(clk), .RN(n3128), .Q(pic_A[12]), 
        .QN(n4724) );
  DFFRX4 \FB_A_reg[1]  ( .D(n1595), .CK(clk), .RN(n3130), .Q(N4410), .QN(n4797) );
  DFFRX4 \offset_reg[13]  ( .D(n1649), .CK(clk), .RN(n3139), .Q(N802), .QN(
        n2989) );
  DFFRX2 \offset_w_reg[8]  ( .D(n1632), .CK(clk), .RN(n3137), .Q(offset_w[8]), 
        .QN(n4729) );
  DFFRX2 \offset_w_reg[1]  ( .D(n1672), .CK(clk), .RN(n3125), .Q(N4346), .QN(
        n4736) );
  DFFRX2 \offset_w_reg[3]  ( .D(n1627), .CK(clk), .RN(n3138), .Q(N4348), .QN(
        n4734) );
  DFFRX2 \offset_w_reg[4]  ( .D(n1628), .CK(clk), .RN(n3137), .Q(N4349), .QN(
        n4733) );
  DFFRX2 \offset_w_reg[5]  ( .D(n1629), .CK(clk), .RN(n3125), .Q(N4350), .QN(
        n4732) );
  DFFRX2 \offset_w_reg[6]  ( .D(n1630), .CK(clk), .RN(n3138), .Q(N4351), .QN(
        n4731) );
  DFFRX4 \offset_reg[12]  ( .D(n1648), .CK(clk), .RN(n3140), .Q(N801), .QN(
        n2990) );
  DFFRX2 \offset_w_reg[13]  ( .D(n1637), .CK(clk), .RN(n3125), .Q(offset_w[13]), .QN(n4739) );
  DFFRX2 \offset_w_reg[11]  ( .D(n1635), .CK(clk), .RN(n3137), .Q(offset_w[11]), .QN(n4741) );
  DFFRX2 \offset_w_reg[2]  ( .D(n1626), .CK(clk), .RN(n3125), .Q(N4347), .QN(
        n4735) );
  DFFRX2 \offset_w_reg[14]  ( .D(n1671), .CK(clk), .RN(n3135), .Q(offset_w[14]), .QN(n4738) );
  DFFRX2 \offset_w_reg[9]  ( .D(n1633), .CK(clk), .RN(n3138), .Q(offset_w[9]), 
        .QN(n4728) );
  DFFRX2 \offset_w_reg[12]  ( .D(n1636), .CK(clk), .RN(n3138), .Q(offset_w[12]), .QN(n4740) );
  DFFRX2 \offset_w_reg[10]  ( .D(n1634), .CK(clk), .RN(n3137), .Q(offset_w[10]), .QN(n4742) );
  DFFRX2 \offset_w_reg[15]  ( .D(n1676), .CK(clk), .RN(n3137), .Q(offset_w[15]), .QN(n4737) );
  DFFRX1 \offset_reg[3]  ( .D(n1640), .CK(clk), .RN(n3135), .QN(n2982) );
  DFFRX4 \offset_reg[14]  ( .D(n1650), .CK(clk), .RN(n3136), .Q(N803), .QN(
        n2985) );
  DFFRX4 \offset_reg[15]  ( .D(n1651), .CK(clk), .RN(n3139), .Q(N804), .QN(
        n2992) );
  DFFRX4 \sec_reg[0]  ( .D(n1625), .CK(clk), .RN(n3141), .Q(N6401), .QN(n4707)
         );
  DFFRX1 \hour_reg[4]  ( .D(hour_n[4]), .CK(clk), .RN(n3125), .Q(hour[4]), 
        .QN(n4861) );
  DFFRX2 \min_reg[3]  ( .D(min_n[3]), .CK(clk), .RN(n3134), .Q(min[3]), .QN(
        n4868) );
  DFFRX2 \min_reg[2]  ( .D(min_n[2]), .CK(clk), .RN(n3136), .Q(N6151), .QN(
        n4867) );
  DFFRX1 \hour_reg[2]  ( .D(hour_n[2]), .CK(clk), .RN(n3131), .Q(hour[2]), 
        .QN(n4863) );
  DFFRX1 \state_reg[0]  ( .D(n1674), .CK(clk), .RN(n3131), .Q(state[0]), .QN(
        n2973) );
  DFFRX2 \pix_c_reg[1]  ( .D(n1678), .CK(clk), .RN(n3127), .QN(n4855) );
  DFFRX2 \hour_reg[0]  ( .D(hour_n[0]), .CK(clk), .RN(n3136), .Q(N5910), .QN(
        n4809) );
  DFFRX1 \min_reg[5]  ( .D(min_n[5]), .CK(clk), .RN(n3125), .Q(min[5]), .QN(
        n4864) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_3  ( .A(N672), .B(N666), .CI(
        \add_0_root_add_0_root_add_209_3/carry[3] ), .CO(
        \add_0_root_add_0_root_add_209_3/carry[4] ), .S(N712) );
  ADDFXL \add_0_root_add_0_root_add_209_3/U1_2  ( .A(N671), .B(n4855), .CI(
        n3102), .CO(\add_0_root_add_0_root_add_209_3/carry[3] ), .S(N711) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_2  ( .A(N1383), .B(n4855), .CI(
        n3103), .CO(\add_0_root_add_1_root_add_282_4/carry[3] ), .S(N1443) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_2  ( .A(N7683), .B(n4855), 
        .CI(n3104), .CO(\add_0_root_add_0_root_add_579_4_cf/carry[3] ), .S(
        N4178) );
  ADDFXL \add_0_root_add_0_root_add_579_4_cf/U1_3  ( .A(N7682), .B(N666), .CI(
        \add_0_root_add_0_root_add_579_4_cf/carry[3] ), .CO(
        \add_0_root_add_0_root_add_579_4_cf/carry[4] ), .S(N4179) );
  ADDFXL \add_0_root_add_0_root_add_446_3/U1_3  ( .A(N2813), .B(N666), .CI(
        \add_0_root_add_0_root_add_446_3/carry[3] ), .CO(
        \add_0_root_add_0_root_add_446_3/carry[4] ), .S(N2853) );
  ADDFXL \add_0_root_add_1_root_add_282_4/U1_3  ( .A(N1384), .B(N666), .CI(
        \add_0_root_add_1_root_add_282_4/carry[3] ), .CO(
        \add_0_root_add_1_root_add_282_4/carry[4] ), .S(N1444) );
  OR2X1 U2444 ( .A(n2953), .B(n3206), .Y(n2952) );
  OA22X1 U2445 ( .A0(n4260), .A1(n3376), .B0(n3244), .B1(n3270), .Y(n2953) );
  AND2X2 U2446 ( .A(n3016), .B(N6160), .Y(n2954) );
  AND2X2 U2447 ( .A(n3016), .B(N6401), .Y(n2955) );
  NOR2X4 U2448 ( .A(pic_size[9]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[9] ), .Y(n2956) );
  XNOR2X1 U2449 ( .A(\gt_332/n15 ), .B(n3305), .Y(N666) );
  CLKINVX1 U2450 ( .A(n3950), .Y(n3946) );
  INVX8 U2451 ( .A(n2982), .Y(n3016) );
  OAI222XL U2452 ( .A0(n3472), .A1(n3767), .B0(n3777), .B1(n3768), .C0(n3770), 
        .C1(n2995), .Y(n1621) );
  AND2X2 U2453 ( .A(n3016), .B(N5910), .Y(n2960) );
  AND2X2 U2454 ( .A(n3015), .B(N7704), .Y(n2962) );
  AND2X1 U2455 ( .A(n4854), .B(n3561), .Y(n2964) );
  AND2X1 U2456 ( .A(n3560), .B(n3306), .Y(n2966) );
  AND2X2 U2457 ( .A(n3015), .B(N2811), .Y(n2969) );
  AND2X2 U2458 ( .A(n3015), .B(N7622), .Y(n2970) );
  AND2X2 U2459 ( .A(n3015), .B(N4325), .Y(n2971) );
  AND2X2 U2460 ( .A(N2422), .B(n3105), .Y(n2972) );
  AND2X2 U2461 ( .A(offset_w[15]), .B(n3086), .Y(n2976) );
  AOI21X4 U2462 ( .A0(n3212), .A1(n3222), .B0(n3195), .Y(n4382) );
  NOR2X2 U2463 ( .A(n3306), .B(n3990), .Y(n3945) );
  INVX3 U2464 ( .A(n4854), .Y(n3306) );
  OAI221X1 U2465 ( .A0(n3450), .A1(n3436), .B0(n3462), .B1(n3463), .C0(n3464), 
        .Y(n3307) );
  OAI211X4 U2466 ( .A0(n3443), .A1(n3316), .B0(n3431), .C0(n3444), .Y(n3189)
         );
  INVX3 U2467 ( .A(IM_Q[9]), .Y(n3470) );
  OAI222XL U2468 ( .A0(n3473), .A1(n3767), .B0(n3768), .B1(n3778), .C0(n3770), 
        .C1(n2994), .Y(n1620) );
  INVX3 U2469 ( .A(IM_Q[1]), .Y(n3473) );
  INVX3 U2470 ( .A(IM_Q[8]), .Y(n3471) );
  INVX3 U2471 ( .A(IM_Q[19]), .Y(n3806) );
  OAI21X1 U2472 ( .A0(n3244), .A1(n3270), .B0(n3284), .Y(n4313) );
  NAND2X2 U2473 ( .A(n3468), .B(n3560), .Y(n3270) );
  OAI211XL U2474 ( .A0(n3270), .A1(n3271), .B0(n3272), .C0(n3273), .Y(n3269)
         );
  OAI211XL U2475 ( .A0(n3270), .A1(n4275), .B0(n4276), .C0(n4277), .Y(n4274)
         );
  INVX3 U2476 ( .A(n3379), .Y(n3449) );
  INVX3 U2477 ( .A(n2964), .Y(n2996) );
  INVX3 U2478 ( .A(IM_Q[2]), .Y(n3472) );
  OAI222XL U2479 ( .A0(n3474), .A1(n3767), .B0(n3768), .B1(n3769), .C0(n3770), 
        .C1(n4707), .Y(n1625) );
  INVX3 U2480 ( .A(IM_Q[0]), .Y(n3474) );
  INVX3 U2481 ( .A(n3944), .Y(n3828) );
  INVX3 U2482 ( .A(n3952), .Y(n3830) );
  INVXL U2483 ( .A(n3225), .Y(n2997) );
  INVX3 U2484 ( .A(n2997), .Y(n2998) );
  NOR2BXL U2485 ( .AN(n3560), .B(n3766), .Y(n3225) );
  OA21X2 U2486 ( .A0(n3181), .A1(n3781), .B0(n3782), .Y(n3770) );
  AOI22XL U2487 ( .A0(N5865), .A1(n3829), .B0(N5968), .B1(n3830), .Y(n3942) );
  AOI22XL U2488 ( .A0(N5864), .A1(n3829), .B0(N5967), .B1(n3830), .Y(n3930) );
  AOI22XL U2489 ( .A0(N5863), .A1(n3829), .B0(N5966), .B1(n3830), .Y(n3918) );
  AOI22XL U2490 ( .A0(N5862), .A1(n3829), .B0(N5965), .B1(n3830), .Y(n3906) );
  AOI22XL U2491 ( .A0(n3074), .A1(n3829), .B0(n3074), .B1(n3830), .Y(n3894) );
  AOI22XL U2492 ( .A0(n3016), .A1(n3829), .B0(n3016), .B1(n3830), .Y(n3882) );
  INVX3 U2493 ( .A(n3953), .Y(n3829) );
  NAND3X2 U2494 ( .A(n3990), .B(n4004), .C(n4202), .Y(n4023) );
  NOR2BX2 U2495 ( .AN(n3560), .B(n3379), .Y(n3237) );
  NAND3X2 U2496 ( .A(n2965), .B(n2958), .C(pic_size[8]), .Y(n3379) );
  OA21X2 U2497 ( .A0(n3987), .A1(n3988), .B0(n3820), .Y(n3819) );
  NOR2X2 U2498 ( .A(n3784), .B(n3354), .Y(n3820) );
  INVXL U2499 ( .A(n4395), .Y(n2999) );
  INVX3 U2500 ( .A(n2999), .Y(n3000) );
  NOR2BXL U2501 ( .AN(n2998), .B(n3436), .Y(n4395) );
  INVX3 U2502 ( .A(n2952), .Y(n3001) );
  INVX3 U2503 ( .A(n2966), .Y(n3002) );
  INVX12 U2504 ( .A(n1412), .Y(CR_A[8]) );
  INVX12 U2505 ( .A(n1413), .Y(CR_A[7]) );
  INVX12 U2506 ( .A(n1414), .Y(CR_A[6]) );
  INVX12 U2507 ( .A(n1415), .Y(CR_A[5]) );
  INVX12 U2508 ( .A(n1416), .Y(CR_A[4]) );
  INVX12 U2509 ( .A(n1417), .Y(CR_A[3]) );
  INVX12 U2510 ( .A(n1418), .Y(CR_A[2]) );
  INVX12 U2511 ( .A(n1419), .Y(CR_A[1]) );
  INVX12 U2512 ( .A(n1420), .Y(CR_A[0]) );
  NOR2X4 U2513 ( .A(n4201), .B(n4024), .Y(n4137) );
  CLKINVX2 U2514 ( .A(n4205), .Y(n4201) );
  NOR3X4 U2515 ( .A(n3202), .B(N2136), .C(n3331), .Y(n4141) );
  NAND2X4 U2516 ( .A(N444), .B(n3367), .Y(n3202) );
  NAND2BX4 U2517 ( .AN(n3990), .B(n3306), .Y(n3348) );
  NOR2BX4 U2518 ( .AN(n3522), .B(n3523), .Y(n3489) );
  INVXL U2519 ( .A(n4305), .Y(n3012) );
  INVX3 U2520 ( .A(n3012), .Y(n3013) );
  NOR2BXL U2521 ( .AN(n3237), .B(n3244), .Y(n4305) );
  AND4X4 U2522 ( .A(n3461), .B(n3642), .C(n3643), .D(n3644), .Y(n3484) );
  NAND2X2 U2523 ( .A(n3560), .B(n3950), .Y(n4024) );
  NOR2X2 U2524 ( .A(n3761), .B(n3950), .Y(n3222) );
  NAND4XL U2525 ( .A(n3950), .B(n3002), .C(n3348), .D(n3528), .Y(n3987) );
  NAND2X4 U2526 ( .A(n4854), .B(n3560), .Y(n3950) );
  OAI211XL U2527 ( .A0(n3484), .A1(n2992), .B0(n3494), .C0(n3495), .Y(n1651)
         );
  NAND2X4 U2528 ( .A(n3997), .B(n3459), .Y(n3992) );
  AND4X4 U2529 ( .A(n3459), .B(n4002), .C(n4003), .D(n3457), .Y(n3991) );
  NOR2XL U2530 ( .A(N804), .B(N803), .Y(n3180) );
  INVX4 U2531 ( .A(n4202), .Y(n3623) );
  NOR2X8 U2532 ( .A(n3305), .B(n4257), .Y(n3560) );
  INVXL U2533 ( .A(N4429), .Y(n3014) );
  INVX8 U2534 ( .A(n3014), .Y(n3015) );
  INVX12 U2535 ( .A(\r1712/carry[4] ), .Y(N668) );
  NAND2BXL U2536 ( .AN(\gt_332/n9 ), .B(n3143), .Y(\r1712/carry[4] ) );
  AOI2BB1X4 U2537 ( .A0N(n3525), .A1N(n3526), .B0(n3447), .Y(n3487) );
  NOR3XL U2538 ( .A(n3379), .B(n3440), .C(n3416), .Y(n3526) );
  NOR2BX4 U2539 ( .AN(n3641), .B(n3421), .Y(n3490) );
  OAI33XL U2540 ( .A0(n3415), .A1(n3592), .A2(n3440), .B0(n3328), .B1(n3342), 
        .B2(n3527), .Y(n3641) );
  INVX12 U2541 ( .A(n3017), .Y(IM_D[9]) );
  INVX12 U2542 ( .A(n3019), .Y(IM_D[10]) );
  INVX12 U2543 ( .A(n3021), .Y(IM_D[11]) );
  INVX12 U2544 ( .A(n3023), .Y(IM_D[12]) );
  INVX12 U2545 ( .A(n3025), .Y(IM_D[13]) );
  INVX12 U2546 ( .A(n3027), .Y(IM_D[14]) );
  INVX12 U2547 ( .A(n3029), .Y(IM_D[15]) );
  INVX12 U2548 ( .A(n3031), .Y(IM_D[16]) );
  INVX12 U2549 ( .A(n3033), .Y(IM_D[17]) );
  INVX12 U2550 ( .A(n3035), .Y(IM_D[18]) );
  INVX12 U2551 ( .A(n3037), .Y(IM_D[19]) );
  INVX12 U2552 ( .A(n3039), .Y(IM_D[20]) );
  INVX12 U2553 ( .A(n3041), .Y(IM_D[21]) );
  INVX12 U2554 ( .A(n3043), .Y(IM_D[22]) );
  INVX12 U2555 ( .A(n3045), .Y(IM_D[23]) );
  AOI222XL U2556 ( .A0(n4141), .A1(IM_Q[23]), .B0(n4142), .B1(n4963), .C0(
        n4143), .C1(\IM_D_t[0][23] ), .Y(n4196) );
  AOI22XL U2557 ( .A0(N3222), .A1(n3490), .B0(n93), .B1(n3491), .Y(n3504) );
  AOI22XL U2558 ( .A0(N3223), .A1(n3490), .B0(n92), .B1(n3491), .Y(n3492) );
  AOI22XL U2559 ( .A0(N3224), .A1(n3490), .B0(n91), .B1(n3491), .Y(n3502) );
  AOI22XL U2560 ( .A0(N3226), .A1(n3490), .B0(n89), .B1(n3491), .Y(n3498) );
  AOI22XL U2561 ( .A0(N3225), .A1(n3490), .B0(n90), .B1(n3491), .Y(n3500) );
  AOI22XL U2562 ( .A0(N3214), .A1(n3490), .B0(n101), .B1(n3491), .Y(n3520) );
  OAI211X4 U2563 ( .A0(n3435), .A1(n3523), .B0(n3529), .C0(n3530), .Y(n3491)
         );
  INVX3 U2564 ( .A(n3955), .Y(n3848) );
  OAI21X4 U2565 ( .A0(n2996), .A1(n4201), .B0(n4034), .Y(n4140) );
  OAI221X4 U2566 ( .A0(n3202), .A1(n3477), .B0(n3950), .B1(n4201), .C0(n4204), 
        .Y(n4143) );
  NOR2BX2 U2567 ( .AN(n3967), .B(n3962), .Y(n3843) );
  NAND4XL U2568 ( .A(offset_w[9]), .B(offset_w[8]), .C(N4352), .D(offset_w[14]), .Y(n3176) );
  NOR3X4 U2569 ( .A(n3440), .B(n3421), .C(n3524), .Y(n3488) );
  NAND4X1 U2570 ( .A(n2967), .B(n2959), .C(n2975), .D(n4624), .Y(n4605) );
  INVX3 U2571 ( .A(n3427), .Y(n3190) );
  AND2X2 U2572 ( .A(n3975), .B(n3976), .Y(n3846) );
  OA22X2 U2573 ( .A0(n3945), .A1(n3990), .B0(n3373), .B1(n4004), .Y(n4027) );
  NOR2X2 U2574 ( .A(n3331), .B(n3202), .Y(n3195) );
  INVX3 U2575 ( .A(n3295), .Y(n3208) );
  NOR2X2 U2576 ( .A(n3963), .B(n3961), .Y(n3839) );
  OAI31X1 U2577 ( .A0(sec[3]), .A1(sec[6]), .A2(sec[4]), .B0(n3964), .Y(n3961)
         );
  NAND4XL U2578 ( .A(offset_w[13]), .B(offset_w[12]), .C(offset_w[11]), .D(
        offset_w[10]), .Y(n3177) );
  INVX4 U2579 ( .A(n4121), .Y(n4016) );
  NAND3XL U2580 ( .A(n3340), .B(n4217), .C(n4218), .Y(n4121) );
  OAI211XL U2581 ( .A0(n3484), .A1(n2990), .B0(n3500), .C0(n3501), .Y(n1648)
         );
  OAI211XL U2582 ( .A0(n3201), .A1(n3202), .B0(n3203), .C0(n3204), .Y(n3196)
         );
  NAND3XL U2583 ( .A(n3661), .B(n3379), .C(n3201), .Y(n3482) );
  INVX3 U2584 ( .A(n4244), .Y(n4036) );
  NAND2XL U2585 ( .A(n3449), .B(n3338), .Y(n3349) );
  INVX3 U2586 ( .A(n3528), .Y(n3338) );
  AND4X2 U2587 ( .A(n4238), .B(n4211), .C(n4239), .D(n4240), .Y(n4029) );
  AOI22XL U2588 ( .A0(N3741), .A1(n4398), .B0(N4463), .B1(n4399), .Y(n4409) );
  AOI22XL U2589 ( .A0(N3742), .A1(n4398), .B0(N4464), .B1(n4399), .Y(n4426) );
  AOI22XL U2590 ( .A0(N3743), .A1(n4398), .B0(N4465), .B1(n4399), .Y(n4443) );
  AOI22XL U2591 ( .A0(N3744), .A1(n4398), .B0(N4466), .B1(n4399), .Y(n4460) );
  AOI22XL U2592 ( .A0(N3745), .A1(n4398), .B0(N4467), .B1(n4399), .Y(n4477) );
  AOI22XL U2593 ( .A0(N3746), .A1(n4398), .B0(N4468), .B1(n4399), .Y(n4494) );
  AOI22XL U2594 ( .A0(N3747), .A1(n4398), .B0(N4469), .B1(n4399), .Y(n4511) );
  AOI22XL U2595 ( .A0(N3748), .A1(n4398), .B0(N4470), .B1(n4399), .Y(n4528) );
  AOI22XL U2596 ( .A0(N3749), .A1(n4398), .B0(N4471), .B1(n4399), .Y(n4545) );
  AOI22XL U2597 ( .A0(N3750), .A1(n4398), .B0(N4472), .B1(n4399), .Y(n4562) );
  AOI22XL U2598 ( .A0(N3751), .A1(n4398), .B0(N4473), .B1(n4399), .Y(n4581) );
  AOI22XL U2599 ( .A0(N3740), .A1(n4398), .B0(N4462), .B1(n4399), .Y(n4386) );
  NOR3BX1 U2600 ( .AN(n3459), .B(n3340), .C(n3367), .Y(n4007) );
  NOR3X2 U2601 ( .A(n3354), .B(n3423), .C(n3206), .Y(n3459) );
  AOI31X4 U2602 ( .A0(n3422), .A1(n3478), .A2(n3764), .B0(n3482), .Y(n3310) );
  NOR2X2 U2603 ( .A(n4605), .B(n3451), .Y(n3422) );
  CLKINVX3 U2604 ( .A(n3371), .Y(n3244) );
  NOR2X2 U2605 ( .A(n3463), .B(n3478), .Y(n3371) );
  NOR2X2 U2606 ( .A(n3761), .B(n3528), .Y(n3218) );
  NAND2X2 U2607 ( .A(n3561), .B(n3306), .Y(n3528) );
  NAND2X2 U2608 ( .A(n4871), .B(n3712), .Y(n3761) );
  INVX3 U2609 ( .A(n3297), .Y(n3241) );
  AO22X2 U2610 ( .A0(n3839), .A1(n3945), .B0(n3338), .B1(n3847), .Y(n3831) );
  NOR2X2 U2611 ( .A(n3975), .B(n3973), .Y(n3847) );
  AO22X2 U2612 ( .A0(n3838), .A1(n3945), .B0(n3338), .B1(n3846), .Y(n3827) );
  NOR2BX2 U2613 ( .AN(n3963), .B(n3961), .Y(n3838) );
  AND2XL U2614 ( .A(offset_w[9]), .B(offset_w[8]), .Y(n3091) );
  NOR2X4 U2615 ( .A(n4201), .B(n4027), .Y(n4133) );
  OAI211XL U2616 ( .A0(n3484), .A1(n2989), .B0(n3498), .C0(n3499), .Y(n1649)
         );
  AND2X2 U2617 ( .A(n4608), .B(n2973), .Y(n3357) );
  INVX3 U2618 ( .A(n4579), .Y(n3219) );
  OA22XL U2619 ( .A0(n3471), .A1(n4656), .B0(n4810), .B1(n4657), .Y(n4643) );
  INVX2 U2620 ( .A(n4639), .Y(n4657) );
  INVX3 U2621 ( .A(n3483), .Y(n4032) );
  INVX3 U2622 ( .A(n3951), .Y(n3852) );
  INVX3 U2623 ( .A(n4605), .Y(n3531) );
  NOR2BX2 U2624 ( .AN(n3561), .B(n3451), .Y(n3235) );
  NAND3X2 U2625 ( .A(n2974), .B(n2958), .C(pic_size[7]), .Y(n3451) );
  NOR3X2 U2626 ( .A(n3426), .B(n1424), .C(n3712), .Y(n3332) );
  NOR3BX1 U2627 ( .AN(n3431), .B(n3340), .C(n3367), .Y(n3475) );
  OAI22X1 U2628 ( .A0(n3369), .A1(n2973), .B0(n4263), .B1(n4264), .Y(n3431) );
  INVX3 U2629 ( .A(n3798), .Y(n3367) );
  MXI2XL U2630 ( .A(n2068), .B(n3993), .S0(n4006), .Y(n1560) );
  MXI2XL U2631 ( .A(n2069), .B(n3994), .S0(n4006), .Y(n1559) );
  MXI2XL U2632 ( .A(n2070), .B(n3995), .S0(n4006), .Y(n1558) );
  MXI2XL U2633 ( .A(n2071), .B(n3996), .S0(n4006), .Y(n1557) );
  MXI2XL U2634 ( .A(n2072), .B(n3806), .S0(n4006), .Y(n1556) );
  MXI2XL U2635 ( .A(n2073), .B(n3808), .S0(n4006), .Y(n1555) );
  MXI2XL U2636 ( .A(n2074), .B(n3809), .S0(n4006), .Y(n1554) );
  MXI2XL U2637 ( .A(n2075), .B(n3810), .S0(n4006), .Y(n1553) );
  MXI2XL U2638 ( .A(n2076), .B(n3811), .S0(n4006), .Y(n1552) );
  MXI2XL U2639 ( .A(n2077), .B(n3812), .S0(n4006), .Y(n1551) );
  MXI2XL U2640 ( .A(n2078), .B(n3813), .S0(n4006), .Y(n1550) );
  MXI2XL U2641 ( .A(n2079), .B(n3814), .S0(n4006), .Y(n1549) );
  MXI2XL U2642 ( .A(n2080), .B(n3815), .S0(n4006), .Y(n1548) );
  MXI2XL U2643 ( .A(n2081), .B(n3816), .S0(n4006), .Y(n1547) );
  MXI2XL U2644 ( .A(n2082), .B(n3470), .S0(n4006), .Y(n1546) );
  MXI2XL U2645 ( .A(n2083), .B(n3471), .S0(n4006), .Y(n1545) );
  MXI2XL U2646 ( .A(n4746), .B(n3299), .S0(n4006), .Y(n1544) );
  MXI2XL U2647 ( .A(n4747), .B(n3779), .S0(n4006), .Y(n1543) );
  MXI2XL U2648 ( .A(n4748), .B(n3771), .S0(n4006), .Y(n1542) );
  MXI2XL U2649 ( .A(n4749), .B(n3773), .S0(n4006), .Y(n1541) );
  MXI2XL U2650 ( .A(n4750), .B(n3775), .S0(n4006), .Y(n1540) );
  MXI2XL U2651 ( .A(n4751), .B(n3472), .S0(n4006), .Y(n1539) );
  MXI2XL U2652 ( .A(n4752), .B(n3473), .S0(n4006), .Y(n1538) );
  MXI2XL U2653 ( .A(n4753), .B(n3474), .S0(n4006), .Y(n1537) );
  INVX3 U2654 ( .A(\sub_609/carry[4] ), .Y(N4433) );
  NAND2BXL U2655 ( .AN(\gt_332/n9 ), .B(n3142), .Y(\sub_609/carry[4] ) );
  NAND2X2 U2656 ( .A(n3372), .B(n3761), .Y(n3347) );
  CLKINVX2 U2657 ( .A(n3451), .Y(n3372) );
  NOR2BX4 U2658 ( .AN(n3226), .B(n3436), .Y(n4393) );
  AOI22XL U2659 ( .A0(N4107), .A1(n2998), .B0(N4365), .B1(n3226), .Y(n3274) );
  AOI22XL U2660 ( .A0(N4106), .A1(n2998), .B0(N4364), .B1(n3226), .Y(n3214) );
  AOI22XL U2661 ( .A0(N4108), .A1(n2998), .B0(N4366), .B1(n3226), .Y(n4618) );
  AOI22XL U2662 ( .A0(N4109), .A1(n2998), .B0(N4367), .B1(n3226), .Y(n4287) );
  AOI22XL U2663 ( .A0(N4113), .A1(n2998), .B0(N4371), .B1(n3226), .Y(n4369) );
  NOR2X2 U2664 ( .A(n4004), .B(n3766), .Y(n3226) );
  NOR2BX2 U2665 ( .AN(n3981), .B(n3974), .Y(n3851) );
  INVX16 U2666 ( .A(n1423), .Y(IM_A[0]) );
  INVX12 U2667 ( .A(n4840), .Y(IM_A[4]) );
  INVX12 U2668 ( .A(n4839), .Y(IM_A[5]) );
  INVX12 U2669 ( .A(n4838), .Y(IM_A[6]) );
  INVX12 U2670 ( .A(n4837), .Y(IM_A[7]) );
  BUFX12 U2671 ( .A(n4962), .Y(IM_A[8]) );
  BUFX12 U2672 ( .A(n4961), .Y(IM_A[9]) );
  BUFX12 U2673 ( .A(n4960), .Y(IM_A[10]) );
  BUFX12 U2674 ( .A(n4959), .Y(IM_A[11]) );
  BUFX12 U2675 ( .A(n4958), .Y(IM_A[12]) );
  BUFX12 U2676 ( .A(n4957), .Y(IM_A[13]) );
  BUFX12 U2677 ( .A(n4956), .Y(IM_A[14]) );
  BUFX12 U2678 ( .A(n4955), .Y(IM_A[15]) );
  BUFX12 U2679 ( .A(n4954), .Y(IM_A[16]) );
  BUFX12 U2680 ( .A(n4953), .Y(IM_A[17]) );
  BUFX12 U2681 ( .A(n4952), .Y(IM_A[18]) );
  BUFX12 U2682 ( .A(n4951), .Y(IM_A[19]) );
  AOI22XL U2683 ( .A0(N3636), .A1(n4396), .B0(N3771), .B1(n4397), .Y(n4582) );
  AOI22XL U2684 ( .A0(N3635), .A1(n4396), .B0(N3770), .B1(n4397), .Y(n4563) );
  AOI22XL U2685 ( .A0(N3634), .A1(n4396), .B0(N3769), .B1(n4397), .Y(n4546) );
  AOI22XL U2686 ( .A0(N3633), .A1(n4396), .B0(N3768), .B1(n4397), .Y(n4529) );
  AOI22XL U2687 ( .A0(N3632), .A1(n4396), .B0(N3767), .B1(n4397), .Y(n4512) );
  AOI22XL U2688 ( .A0(N3631), .A1(n4396), .B0(N3766), .B1(n4397), .Y(n4495) );
  NOR2BX2 U2689 ( .AN(n3218), .B(n3436), .Y(n4397) );
  AOI22XL U2690 ( .A0(N3625), .A1(n4396), .B0(N3760), .B1(n4397), .Y(n4387) );
  AOI22XL U2691 ( .A0(N3626), .A1(n4396), .B0(N3761), .B1(n4397), .Y(n4410) );
  AOI22XL U2692 ( .A0(N3627), .A1(n4396), .B0(N3762), .B1(n4397), .Y(n4427) );
  AOI22XL U2693 ( .A0(N3628), .A1(n4396), .B0(N3763), .B1(n4397), .Y(n4444) );
  AOI22XL U2694 ( .A0(N3629), .A1(n4396), .B0(N3764), .B1(n4397), .Y(n4461) );
  AOI22XL U2695 ( .A0(N3630), .A1(n4396), .B0(N3765), .B1(n4397), .Y(n4478) );
  AND4X4 U2696 ( .A(n3522), .B(n3661), .C(n3422), .D(n3478), .Y(n3312) );
  NOR2BX4 U2697 ( .AN(n4200), .B(n3202), .Y(n4134) );
  MXI2XL U2698 ( .A(n4789), .B(n3470), .S0(n3807), .Y(n1603) );
  OAI211XL U2699 ( .A0(n3484), .A1(n2988), .B0(n3502), .C0(n3503), .Y(n1647)
         );
  INVX3 U2700 ( .A(n3415), .Y(n3343) );
  AOI2BB1X2 U2701 ( .A0N(n3410), .A1N(n3433), .B0(n3415), .Y(n4014) );
  NAND3X2 U2702 ( .A(n2965), .B(n2974), .C(pic_size[9]), .Y(n3415) );
  INVX3 U2703 ( .A(n3954), .Y(n3840) );
  OAI22X2 U2704 ( .A0(n3954), .A1(n3949), .B0(n3528), .B1(n3955), .Y(n3832) );
  OAI222X4 U2705 ( .A0(n3528), .A1(n3947), .B0(n3948), .B1(n3949), .C0(n3950), 
        .C1(n3951), .Y(n3826) );
  CLKINVX2 U2706 ( .A(n3945), .Y(n3949) );
  MXI2XL U2707 ( .A(n4708), .B(n3470), .S0(n4262), .Y(n1453) );
  MXI2XL U2708 ( .A(n4709), .B(n3471), .S0(n4262), .Y(n1452) );
  NOR3BX1 U2709 ( .AN(n3787), .B(n3788), .C(n4874), .Y(n3353) );
  NOR2X2 U2710 ( .A(n3188), .B(N6483), .Y(n3787) );
  INVX3 U2711 ( .A(N444), .Y(n3478) );
  NOR2X2 U2712 ( .A(n3463), .B(N444), .Y(n3210) );
  OAI211XL U2713 ( .A0(N444), .A1(n3375), .B0(n3379), .C0(n3377), .Y(n3466) );
  AOI2BB1X2 U2714 ( .A0N(n3175), .A1N(n3174), .B0(n3173), .Y(N444) );
  INVX3 U2715 ( .A(\sub_601/carry[4] ), .Y(N4323) );
  NOR2X2 U2716 ( .A(n3854), .B(n3852), .Y(n3853) );
  NAND3X2 U2717 ( .A(n4860), .B(n3985), .C(n4859), .Y(n3854) );
  MXI2XL U2718 ( .A(n2975), .B(n3474), .S0(n3300), .Y(n1655) );
  MXI2XL U2719 ( .A(n2967), .B(n3473), .S0(n3300), .Y(n1656) );
  MXI2XL U2720 ( .A(n2959), .B(n3472), .S0(n3300), .Y(n1657) );
  MXI2XL U2721 ( .A(n2974), .B(n3471), .S0(n3300), .Y(n1662) );
  MXI2XL U2722 ( .A(n2958), .B(n3470), .S0(n3300), .Y(n1663) );
  AND3X2 U2723 ( .A(n3475), .B(n3476), .C(n3364), .Y(n3300) );
  NOR2BX4 U2724 ( .AN(n3224), .B(n3436), .Y(n4394) );
  NOR2BX2 U2725 ( .AN(n3561), .B(n3766), .Y(n3224) );
  INVX3 U2726 ( .A(n3316), .Y(n3410) );
  NOR2XL U2727 ( .A(n3347), .B(n3316), .Y(n4205) );
  OAI211X4 U2728 ( .A0(n4206), .A1(n3316), .B0(n4207), .C0(n4208), .Y(n4142)
         );
  OAI32X4 U2729 ( .A0(n3417), .A1(n4202), .A2(n3202), .B0(n3316), .B1(n4203), 
        .Y(n4135) );
  NAND2X2 U2730 ( .A(n3360), .B(n3531), .Y(n3316) );
  INVX3 U2731 ( .A(n4203), .Y(n4018) );
  NAND2XL U2732 ( .A(n3449), .B(n3623), .Y(n4203) );
  NOR2X2 U2733 ( .A(n3981), .B(n3849), .Y(n3850) );
  INVX3 U2734 ( .A(n3947), .Y(n3849) );
  MXI2XL U2735 ( .A(n4798), .B(n3806), .S0(n3807), .Y(n1613) );
  NAND2X2 U2736 ( .A(n3781), .B(n3354), .Y(n4656) );
  CLKINVX2 U2737 ( .A(n3199), .Y(n3354) );
  NOR2BX4 U2738 ( .AN(n3238), .B(n3244), .Y(n4304) );
  NOR2BX2 U2739 ( .AN(n3561), .B(n3379), .Y(n3238) );
  AO22XL U2740 ( .A0(N808), .A1(n3239), .B0(N710), .B1(n3238), .Y(n3281) );
  NAND2XL U2741 ( .A(N1442), .B(n3238), .Y(n3272) );
  NAND2XL U2742 ( .A(N712), .B(n3238), .Y(n4276) );
  AOI22XL U2743 ( .A0(N1441), .A1(n3238), .B0(n3239), .B1(N944), .Y(n3227) );
  NOR2BX4 U2744 ( .AN(n3221), .B(n3436), .Y(n4398) );
  NOR2X2 U2745 ( .A(n2996), .B(n3761), .Y(n3221) );
  NOR2BX4 U2746 ( .AN(n3220), .B(n3436), .Y(n4396) );
  NOR2X2 U2747 ( .A(n3761), .B(n3002), .Y(n3220) );
  NAND2X4 U2748 ( .A(n3410), .B(n3372), .Y(n3436) );
  NOR2BX4 U2749 ( .AN(n4028), .B(n4201), .Y(n4136) );
  NOR2BX2 U2750 ( .AN(n3561), .B(n2964), .Y(n4028) );
  NOR2BX4 U2751 ( .AN(n3257), .B(n3244), .Y(n4302) );
  CLKAND2X3 U2752 ( .A(n4217), .B(n3340), .Y(n3240) );
  NAND2XL U2753 ( .A(n3788), .B(n4625), .Y(n4217) );
  INVX2 U2754 ( .A(n3457), .Y(n3340) );
  OAI211XL U2755 ( .A0(n3484), .A1(n2987), .B0(n3492), .C0(n3493), .Y(n1652)
         );
  BUFX4 U2756 ( .A(n4008), .Y(n3059) );
  MXI2XL U2757 ( .A(n4777), .B(n3474), .S0(n3059), .Y(n1513) );
  MXI2XL U2758 ( .A(n4766), .B(n3473), .S0(n3059), .Y(n1514) );
  MXI2XL U2759 ( .A(n4761), .B(n3472), .S0(n3059), .Y(n1515) );
  MXI2XL U2760 ( .A(n4760), .B(n3775), .S0(n3059), .Y(n1516) );
  MXI2XL U2761 ( .A(n4759), .B(n3773), .S0(n3059), .Y(n1517) );
  MXI2XL U2762 ( .A(n4758), .B(n3771), .S0(n3059), .Y(n1518) );
  NOR2BXL U2763 ( .AN(n4007), .B(n3528), .Y(n4008) );
  MXI2XL U2764 ( .A(n4762), .B(n3993), .S0(n3059), .Y(n1536) );
  MXI2XL U2765 ( .A(n4763), .B(n3994), .S0(n3059), .Y(n1535) );
  MXI2XL U2766 ( .A(n4764), .B(n3995), .S0(n3059), .Y(n1534) );
  MXI2XL U2767 ( .A(n4765), .B(n3996), .S0(n3059), .Y(n1533) );
  MXI2XL U2768 ( .A(n4767), .B(n3806), .S0(n3059), .Y(n1532) );
  MXI2XL U2769 ( .A(n4768), .B(n3808), .S0(n3059), .Y(n1531) );
  MXI2XL U2770 ( .A(n4769), .B(n3809), .S0(n3059), .Y(n1530) );
  MXI2XL U2771 ( .A(n4770), .B(n3810), .S0(n3059), .Y(n1529) );
  MXI2XL U2772 ( .A(n4771), .B(n3811), .S0(n3059), .Y(n1528) );
  MXI2XL U2773 ( .A(n4772), .B(n3812), .S0(n3059), .Y(n1527) );
  MXI2XL U2774 ( .A(n4773), .B(n3813), .S0(n3059), .Y(n1526) );
  MXI2XL U2775 ( .A(n4774), .B(n3814), .S0(n3059), .Y(n1525) );
  MXI2XL U2776 ( .A(n4775), .B(n3815), .S0(n3059), .Y(n1524) );
  MXI2XL U2777 ( .A(n4776), .B(n3816), .S0(n3059), .Y(n1523) );
  MXI2XL U2778 ( .A(n4754), .B(n3470), .S0(n3059), .Y(n1522) );
  MXI2XL U2779 ( .A(n4755), .B(n3471), .S0(n3059), .Y(n1521) );
  MXI2XL U2780 ( .A(n4756), .B(n3299), .S0(n3059), .Y(n1520) );
  MXI2XL U2781 ( .A(n4757), .B(n3779), .S0(n3059), .Y(n1519) );
  NOR2X8 U2782 ( .A(n4257), .B(n4855), .Y(n3561) );
  NAND2X4 U2783 ( .A(n3319), .B(n3531), .Y(n3440) );
  NAND2BX4 U2784 ( .AN(n3328), .B(n3319), .Y(n3248) );
  NAND2X4 U2785 ( .A(n3336), .B(n3319), .Y(n3246) );
  INVX3 U2786 ( .A(n3202), .Y(n3319) );
  OAI21X4 U2787 ( .A0(n3376), .A1(n4580), .B0(n3293), .Y(n4314) );
  OAI21X4 U2788 ( .A0(n3270), .A1(n3376), .B0(n3286), .Y(n4308) );
  NOR2BX4 U2789 ( .AN(n3238), .B(n3376), .Y(n4306) );
  NOR2BX4 U2790 ( .AN(n3235), .B(n3376), .Y(n4303) );
  NOR2BX4 U2791 ( .AN(n3237), .B(n3376), .Y(n4301) );
  CLKINVX3 U2792 ( .A(n3210), .Y(n3376) );
  OAI22X4 U2793 ( .A0(n3244), .A1(n3259), .B0(n3258), .B1(n3376), .Y(n3291) );
  OAI22X4 U2794 ( .A0(n3244), .A1(n3258), .B0(n3259), .B1(n3376), .Y(n3292) );
  AOI2BB1XL U2795 ( .A0N(n3404), .A1N(n3405), .B0(n3316), .Y(n3403) );
  NAND3X2 U2796 ( .A(n2966), .B(n3410), .C(n3405), .Y(n4034) );
  NAND3XL U2797 ( .A(n3410), .B(n3946), .C(n3405), .Y(n4204) );
  NAND3X2 U2798 ( .A(n2964), .B(n3410), .C(n3405), .Y(n4035) );
  NAND2XL U2799 ( .A(n3405), .B(n4257), .Y(n4241) );
  NOR2X2 U2800 ( .A(n3761), .B(n3451), .Y(n3405) );
  OAI21X1 U2801 ( .A0(n4644), .A1(n4645), .B0(n3181), .Y(n4638) );
  NAND3BX2 U2802 ( .AN(n4645), .B(n3181), .C(n4644), .Y(n4626) );
  NAND3BX2 U2803 ( .AN(n4669), .B(n3181), .C(n4645), .Y(n4646) );
  MXI2X2 U2804 ( .A(n4672), .B(n4673), .S0(n4644), .Y(n4645) );
  NOR2BX2 U2805 ( .AN(n3223), .B(n3436), .Y(n4399) );
  AOI22XL U2806 ( .A0(N4455), .A1(n3223), .B0(N4177), .B1(n3224), .Y(n3275) );
  AOI22XL U2807 ( .A0(N4454), .A1(n3223), .B0(N4176), .B1(n3224), .Y(n3215) );
  AOI22XL U2808 ( .A0(N4456), .A1(n3223), .B0(N4178), .B1(n3224), .Y(n4619) );
  AOI22XL U2809 ( .A0(N4461), .A1(n3223), .B0(N4183), .B1(n3224), .Y(n4370) );
  AOI22XL U2810 ( .A0(N4460), .A1(n3223), .B0(N4182), .B1(n3224), .Y(n4352) );
  NOR2X2 U2811 ( .A(n3990), .B(n3766), .Y(n3223) );
  NOR2X2 U2812 ( .A(n3967), .B(n3841), .Y(n3842) );
  INVX3 U2813 ( .A(n3948), .Y(n3841) );
  NAND4BXL U2814 ( .AN(n3260), .B(n3261), .C(n3262), .D(n3263), .Y(n1683) );
  INVX12 U2815 ( .A(n4843), .Y(IM_A[1]) );
  BUFX12 U2816 ( .A(n4985), .Y(IM_D[1]) );
  BUFX12 U2817 ( .A(n4984), .Y(IM_D[2]) );
  BUFX12 U2818 ( .A(n4983), .Y(IM_D[3]) );
  BUFX12 U2819 ( .A(n4982), .Y(IM_D[4]) );
  BUFX12 U2820 ( .A(n4981), .Y(IM_D[5]) );
  BUFX12 U2821 ( .A(n4980), .Y(IM_D[6]) );
  BUFX12 U2822 ( .A(n4979), .Y(IM_D[7]) );
  BUFX12 U2823 ( .A(n4978), .Y(IM_D[8]) );
  BUFX12 U2824 ( .A(n4986), .Y(IM_D[0]) );
  NAND4XL U2825 ( .A(n4265), .B(n4266), .C(n4267), .D(n4268), .Y(n1443) );
  INVX12 U2826 ( .A(n4841), .Y(IM_A[3]) );
  INVX12 U2827 ( .A(n4842), .Y(IM_A[2]) );
  INVX16 U2828 ( .A(n2098), .Y(IM_WEN) );
  XNOR2X1 U2829 ( .A(\gt_332/n9 ), .B(\r1712/carry[3] ), .Y(N667) );
  OAI21X4 U2830 ( .A0(n3467), .A1(n4201), .B0(n4035), .Y(n4138) );
  NOR2BX4 U2831 ( .AN(n4007), .B(n3467), .Y(n4006) );
  AOI32XL U2832 ( .A0(n3372), .A1(n2996), .A2(N444), .B0(n3466), .B1(n3467), 
        .Y(n3462) );
  NAND3XL U2833 ( .A(n3949), .B(n3467), .C(n3952), .Y(n3988) );
  INVX4 U2834 ( .A(n3373), .Y(n3467) );
  OAI21X2 U2835 ( .A0(n3441), .A1(n3442), .B0(n3524), .Y(n4031) );
  OA21X2 U2836 ( .A0(n3436), .A1(n4579), .B0(n3290), .Y(n4381) );
  AND2X2 U2837 ( .A(n4606), .B(n4607), .Y(n3290) );
  XOR2XL U2838 ( .A(N6392), .B(N6391), .Y(N6365) );
  XNOR2XL U2839 ( .A(N6392), .B(N6391), .Y(N6311) );
  AOI22XL U2840 ( .A0(N526), .A1(n4300), .B0(N566), .B1(n4302), .Y(n4567) );
  AOI22XL U2841 ( .A0(N525), .A1(n4300), .B0(N565), .B1(n4302), .Y(n4550) );
  AOI22XL U2842 ( .A0(N524), .A1(n4300), .B0(N564), .B1(n4302), .Y(n4533) );
  AOI22XL U2843 ( .A0(N523), .A1(n4300), .B0(N563), .B1(n4302), .Y(n4516) );
  AOI22XL U2844 ( .A0(N522), .A1(n4300), .B0(N562), .B1(n4302), .Y(n4499) );
  AOI22XL U2845 ( .A0(N521), .A1(n4300), .B0(N561), .B1(n4302), .Y(n4482) );
  NOR2BX4 U2846 ( .AN(n3254), .B(n3244), .Y(n4300) );
  AOI22XL U2847 ( .A0(N4633), .A1(n3312), .B0(n84), .B1(n3313), .Y(n3659) );
  AOI22XL U2848 ( .A0(N4634), .A1(n3312), .B0(n83), .B1(n3313), .Y(n3658) );
  AOI22XL U2849 ( .A0(N4635), .A1(n3312), .B0(n82), .B1(n3313), .Y(n3657) );
  AOI22XL U2850 ( .A0(N4636), .A1(n3312), .B0(n81), .B1(n3313), .Y(n3656) );
  AOI22XL U2851 ( .A0(N4637), .A1(n3312), .B0(n80), .B1(n3313), .Y(n3655) );
  AOI22XL U2852 ( .A0(N4638), .A1(n3312), .B0(n79), .B1(n3313), .Y(n3654) );
  NOR2BX4 U2853 ( .AN(n3660), .B(n3479), .Y(n3313) );
  MXI2XL U2854 ( .A(n4808), .B(n3474), .S0(n3807), .Y(n1594) );
  MXI2XL U2855 ( .A(n4797), .B(n3473), .S0(n3807), .Y(n1595) );
  MXI2XL U2856 ( .A(n4796), .B(n3472), .S0(n3807), .Y(n1596) );
  AND2X4 U2857 ( .A(n3786), .B(n3364), .Y(n3807) );
  MXI2XL U2858 ( .A(n4727), .B(n3474), .S0(n4262), .Y(n1444) );
  MXI2XL U2859 ( .A(n4716), .B(n3473), .S0(n4262), .Y(n1445) );
  MXI2XL U2860 ( .A(n4715), .B(n3472), .S0(n4262), .Y(n1446) );
  MXI2XL U2861 ( .A(n4714), .B(n3775), .S0(n4262), .Y(n1447) );
  MXI2XL U2862 ( .A(n4713), .B(n3773), .S0(n4262), .Y(n1448) );
  MXI2XL U2863 ( .A(n4712), .B(n3771), .S0(n4262), .Y(n1449) );
  AND3X4 U2864 ( .A(n3475), .B(n3476), .C(n3781), .Y(n4262) );
  MXI2XL U2865 ( .A(n4799), .B(n3808), .S0(n3807), .Y(n1612) );
  NOR2X4 U2866 ( .A(n3665), .B(n3202), .Y(n3243) );
  INVX3 U2867 ( .A(n3187), .Y(n3181) );
  AOI2BB1X2 U2868 ( .A0N(n4645), .A1N(n4669), .B0(n3187), .Y(n4648) );
  NAND4X4 U2869 ( .A(n4685), .B(n4686), .C(n4687), .D(n4688), .Y(n3187) );
  CLKBUFX6 U2870 ( .A(n1927), .Y(n3069) );
  CLKINVX4 U2871 ( .A(n1927), .Y(n3381) );
  NAND2XL U2872 ( .A(n3343), .B(n3069), .Y(n3383) );
  MXI2XL U2873 ( .A(N3737), .B(N2323), .S0(n3069), .Y(n3679) );
  MXI2XL U2874 ( .A(N2420), .B(N2334), .S0(n3069), .Y(n3680) );
  MXI2XL U2875 ( .A(N3738), .B(N2324), .S0(n3069), .Y(n3688) );
  MXI2XL U2876 ( .A(N2419), .B(N2333), .S0(n3069), .Y(n3699) );
  OAI211XL U2877 ( .A0(n3484), .A1(n2986), .B0(n3504), .C0(n3505), .Y(n1646)
         );
  OAI21X4 U2878 ( .A0(n3949), .A1(n4201), .B0(n4033), .Y(n4139) );
  NAND3X2 U2879 ( .A(n3338), .B(n3410), .C(n3405), .Y(n4033) );
  BUFX4 U2880 ( .A(n4009), .Y(n3070) );
  INVX8 U2881 ( .A(n4855), .Y(n3305) );
  CLKBUFX8 U2882 ( .A(N791), .Y(n3071) );
  CLKBUFX8 U2883 ( .A(N790), .Y(n3072) );
  CLKBUFX8 U2884 ( .A(N797), .Y(n3073) );
  INVX8 U2885 ( .A(n3074), .Y(n3075) );
  INVX8 U2886 ( .A(n3076), .Y(n3077) );
  INVX8 U2887 ( .A(n3078), .Y(n3079) );
  INVX8 U2888 ( .A(n3080), .Y(n3081) );
  INVX8 U2889 ( .A(n3082), .Y(n3083) );
  CLKINVX1 U2890 ( .A(\r1712/carry[3] ), .Y(n3143) );
  OR2X1 U2891 ( .A(\gt_332/n9 ), .B(\gt_332/n15 ), .Y(\sub_601/carry[4] ) );
  CLKINVX1 U2892 ( .A(n3097), .Y(n3142) );
  XOR2X1 U2893 ( .A(n3073), .B(n3116), .Y(N5856) );
  XOR2X1 U2894 ( .A(n3073), .B(n3117), .Y(N6019) );
  OR2X1 U2895 ( .A(pic_size[2]), .B(pic_size[1]), .Y(
        \sub_2_root_sub_0_root_add_266_3/carry[3] ) );
  OR2X1 U2896 ( .A(N6392), .B(N6391), .Y(\sub_819/carry[3] ) );
  AND2X2 U2897 ( .A(N6392), .B(N6391), .Y(n3084) );
  OR2X1 U2898 ( .A(N6392), .B(N6391), .Y(\sub_827/carry[3] ) );
  OR2X1 U2899 ( .A(N6151), .B(N6150), .Y(\sub_791/carry[3] ) );
  AND2X2 U2900 ( .A(N6151), .B(N6150), .Y(n3085) );
  OR2X1 U2901 ( .A(N6151), .B(N6150), .Y(\sub_799/carry[3] ) );
  OR2X1 U2902 ( .A(hour[2]), .B(N5926), .Y(\sub_767/carry[3] ) );
  AND2X2 U2903 ( .A(offset_w[14]), .B(n3087), .Y(n3086) );
  AND2X2 U2904 ( .A(offset_w[13]), .B(n3088), .Y(n3087) );
  AND2X2 U2905 ( .A(offset_w[12]), .B(n3089), .Y(n3088) );
  AND2X2 U2906 ( .A(offset_w[11]), .B(n3090), .Y(n3089) );
  AND2X2 U2907 ( .A(offset_w[10]), .B(n3091), .Y(n3090) );
  OR2X1 U2908 ( .A(pic_size[8]), .B(\sub_2_root_sub_0_root_add_266_3/carry[8] ), .Y(\sub_2_root_sub_0_root_add_266_3/carry[9] ) );
  OR2X1 U2909 ( .A(pic_size[7]), .B(\sub_2_root_sub_0_root_add_266_3/carry[7] ), .Y(\sub_2_root_sub_0_root_add_266_3/carry[8] ) );
  OR2X1 U2910 ( .A(pic_size[6]), .B(\sub_2_root_sub_0_root_add_266_3/carry[6] ), .Y(\sub_2_root_sub_0_root_add_266_3/carry[7] ) );
  OR2X1 U2911 ( .A(pic_size[5]), .B(\sub_2_root_sub_0_root_add_266_3/carry[5] ), .Y(\sub_2_root_sub_0_root_add_266_3/carry[6] ) );
  OR2X1 U2912 ( .A(pic_size[4]), .B(\sub_2_root_sub_0_root_add_266_3/carry[4] ), .Y(\sub_2_root_sub_0_root_add_266_3/carry[5] ) );
  OR2X1 U2913 ( .A(pic_size[3]), .B(\sub_2_root_sub_0_root_add_266_3/carry[3] ), .Y(\sub_2_root_sub_0_root_add_266_3/carry[4] ) );
  XNOR2X1 U2914 ( .A(pic_size[3]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[3] ), .Y(N1242) );
  OR2X1 U2915 ( .A(sec[3]), .B(\sub_827/carry[3] ), .Y(\sub_827/carry[4] ) );
  OR2X1 U2916 ( .A(sec[3]), .B(N6392), .Y(\sub_821/carry[4] ) );
  AND2X2 U2917 ( .A(sec[3]), .B(\sub_819/carry[3] ), .Y(n3092) );
  AND2X2 U2918 ( .A(sec[3]), .B(n3084), .Y(n3093) );
  OR2X1 U2919 ( .A(min[3]), .B(\sub_799/carry[3] ), .Y(\sub_799/carry[4] ) );
  OR2X1 U2920 ( .A(min[3]), .B(N6151), .Y(\sub_793/carry[4] ) );
  AND2X2 U2921 ( .A(min[3]), .B(\sub_791/carry[3] ), .Y(n3094) );
  AND2X2 U2922 ( .A(min[3]), .B(n3085), .Y(n3095) );
  OR2X1 U2923 ( .A(hour[3]), .B(hour[2]), .Y(\sub_769/carry[4] ) );
  AND2X2 U2924 ( .A(hour[3]), .B(\sub_767/carry[3] ), .Y(n3096) );
  XNOR2X1 U2925 ( .A(sec[3]), .B(N6392), .Y(N6339) );
  XOR2X1 U2926 ( .A(sec[3]), .B(\sub_819/carry[3] ), .Y(N6312) );
  XOR2X1 U2927 ( .A(sec[3]), .B(n3084), .Y(N6366) );
  XNOR2X1 U2928 ( .A(N6392), .B(N6391), .Y(N6418) );
  XNOR2X1 U2929 ( .A(sec[3]), .B(\sub_827/carry[3] ), .Y(N6419) );
  XNOR2X1 U2930 ( .A(min[3]), .B(N6151), .Y(N6098) );
  XNOR2X1 U2931 ( .A(N6151), .B(N6150), .Y(N6070) );
  XOR2X1 U2932 ( .A(min[3]), .B(\sub_791/carry[3] ), .Y(N6071) );
  XOR2X1 U2933 ( .A(N6151), .B(N6150), .Y(N6124) );
  XOR2X1 U2934 ( .A(min[3]), .B(n3085), .Y(N6125) );
  XNOR2X1 U2935 ( .A(N6151), .B(N6150), .Y(N6177) );
  XNOR2X1 U2936 ( .A(min[3]), .B(\sub_799/carry[3] ), .Y(N6178) );
  XNOR2X1 U2937 ( .A(hour[3]), .B(hour[2]), .Y(N5928) );
  XOR2X1 U2938 ( .A(hour[3]), .B(\sub_767/carry[3] ), .Y(N5902) );
  XNOR2X1 U2939 ( .A(hour[2]), .B(N5926), .Y(N5901) );
  XNOR2XL U2940 ( .A(pic_size[2]), .B(pic_size[1]), .Y(N1241) );
  OR2X1 U2941 ( .A(\gt_332/n15 ), .B(n3305), .Y(\r1712/carry[3] ) );
  XOR2XL U2942 ( .A(offset_w[15]), .B(n3086), .Y(N4360) );
  XOR2XL U2943 ( .A(offset_w[14]), .B(n3087), .Y(N4359) );
  XOR2XL U2944 ( .A(offset_w[13]), .B(n3088), .Y(N4358) );
  XOR2XL U2945 ( .A(offset_w[12]), .B(n3089), .Y(N4357) );
  XOR2XL U2946 ( .A(offset_w[11]), .B(n3090), .Y(N4356) );
  XOR2XL U2947 ( .A(offset_w[10]), .B(n3091), .Y(N4355) );
  XOR2XL U2948 ( .A(offset_w[9]), .B(offset_w[8]), .Y(N4354) );
  XNOR2X1 U2949 ( .A(pic_size[9]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[9] ), .Y(N1248) );
  XNOR2X1 U2950 ( .A(pic_size[8]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[8] ), .Y(N1247) );
  XNOR2X1 U2951 ( .A(pic_size[7]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[7] ), .Y(N1246) );
  XNOR2X1 U2952 ( .A(pic_size[6]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[6] ), .Y(N1245) );
  XNOR2X1 U2953 ( .A(pic_size[5]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[5] ), .Y(N1244) );
  AND2X2 U2954 ( .A(\gt_332/n15 ), .B(n3305), .Y(n3097) );
  XNOR2XL U2955 ( .A(pic_size[4]), .B(
        \sub_2_root_sub_0_root_add_266_3/carry[4] ), .Y(N1243) );
  NAND2XL U2956 ( .A(sec[4]), .B(\sub_827/carry[4] ), .Y(n3157) );
  XOR2X1 U2957 ( .A(sec[4]), .B(\sub_827/carry[4] ), .Y(N6420) );
  AND2X2 U2958 ( .A(sec[4]), .B(\sub_821/carry[4] ), .Y(n3098) );
  XOR2X1 U2959 ( .A(sec[4]), .B(\sub_821/carry[4] ), .Y(N6340) );
  OR2X1 U2960 ( .A(sec[4]), .B(n3092), .Y(\sub_819/carry[5] ) );
  XNOR2X1 U2961 ( .A(sec[4]), .B(n3092), .Y(N6313) );
  AND2X2 U2962 ( .A(sec[4]), .B(n3093), .Y(n3099) );
  XOR2X1 U2963 ( .A(sec[4]), .B(n3093), .Y(N6367) );
  OR2X1 U2964 ( .A(sec[4]), .B(sec[3]), .Y(\sub_825/carry[5] ) );
  XNOR2X1 U2965 ( .A(sec[4]), .B(sec[3]), .Y(N6394) );
  NAND2X1 U2966 ( .A(min[4]), .B(\sub_799/carry[4] ), .Y(n3145) );
  XOR2X1 U2967 ( .A(min[4]), .B(\sub_799/carry[4] ), .Y(N6179) );
  AND2X2 U2968 ( .A(min[4]), .B(\sub_793/carry[4] ), .Y(n3100) );
  XOR2X1 U2969 ( .A(min[4]), .B(\sub_793/carry[4] ), .Y(N6099) );
  OR2X1 U2970 ( .A(min[4]), .B(n3094), .Y(\sub_791/carry[5] ) );
  XNOR2X1 U2971 ( .A(min[4]), .B(n3094), .Y(N6072) );
  AND2X2 U2972 ( .A(min[4]), .B(n3095), .Y(n3101) );
  XOR2X1 U2973 ( .A(min[4]), .B(n3095), .Y(N6126) );
  OR2X1 U2974 ( .A(min[4]), .B(min[3]), .Y(\sub_797/carry[5] ) );
  XNOR2X1 U2975 ( .A(min[4]), .B(min[3]), .Y(N6153) );
  NAND2X1 U2976 ( .A(hour[4]), .B(\sub_769/carry[4] ), .Y(n3153) );
  XOR2X1 U2977 ( .A(hour[4]), .B(\sub_769/carry[4] ), .Y(N5929) );
  CLKINVX1 U2978 ( .A(n3096), .Y(n3151) );
  XNOR2X1 U2979 ( .A(hour[4]), .B(n3096), .Y(N5903) );
  AND2X2 U2980 ( .A(n3015), .B(N670), .Y(n3102) );
  AND2X2 U2981 ( .A(n3015), .B(N1382), .Y(n3103) );
  AND2X2 U2982 ( .A(n3015), .B(N7684), .Y(n3104) );
  AND2X2 U2983 ( .A(N2421), .B(n3106), .Y(n3105) );
  AND2X2 U2984 ( .A(N2420), .B(n3107), .Y(n3106) );
  AND2X2 U2985 ( .A(N2419), .B(n3108), .Y(n3107) );
  AND2X2 U2986 ( .A(N2418), .B(n3109), .Y(n3108) );
  AND2X2 U2987 ( .A(N2417), .B(n3110), .Y(n3109) );
  AND2X2 U2988 ( .A(N2416), .B(n3111), .Y(n3110) );
  AND2X2 U2989 ( .A(N2415), .B(n3112), .Y(n3111) );
  AND2X2 U2990 ( .A(N2414), .B(N2413), .Y(n3112) );
  OR2X1 U2991 ( .A(count[7]), .B(n3113), .Y(N6490) );
  AND2X2 U2992 ( .A(count[6]), .B(n3114), .Y(n3113) );
  AND2X2 U2993 ( .A(count[5]), .B(\add_3_root_add_0_root_add_869_4/carry[5] ), 
        .Y(n3114) );
  OR2X1 U2994 ( .A(count[4]), .B(count[3]), .Y(
        \add_3_root_add_0_root_add_869_4/carry[5] ) );
  XNOR2XL U2995 ( .A(\gt_332/n9 ), .B(\gt_332/n15 ), .Y(N4322) );
  XNOR2XL U2996 ( .A(\gt_332/n9 ), .B(n3097), .Y(N4432) );
  XOR2XL U2997 ( .A(\gt_332/n15 ), .B(n3305), .Y(N4431) );
  MX4XL U2998 ( .A(\IM_D_t[0][0] ), .B(\IM_D_t[1][0] ), .C(\IM_D_t[2][0] ), 
        .D(\IM_D_t[3][0] ), .S0(n3015), .S1(n3305), .Y(N251) );
  MX4XL U2999 ( .A(\IM_D_t[0][8] ), .B(\IM_D_t[1][8] ), .C(\IM_D_t[2][8] ), 
        .D(\IM_D_t[3][8] ), .S0(n3015), .S1(n3305), .Y(N243) );
  MX4XL U3000 ( .A(\IM_D_t[0][7] ), .B(\IM_D_t[1][7] ), .C(\IM_D_t[2][7] ), 
        .D(\IM_D_t[3][7] ), .S0(n3015), .S1(n3305), .Y(N244) );
  MX4XL U3001 ( .A(\IM_D_t[0][6] ), .B(\IM_D_t[1][6] ), .C(\IM_D_t[2][6] ), 
        .D(\IM_D_t[3][6] ), .S0(n3015), .S1(n3305), .Y(N245) );
  MX4XL U3002 ( .A(\IM_D_t[0][5] ), .B(\IM_D_t[1][5] ), .C(\IM_D_t[2][5] ), 
        .D(\IM_D_t[3][5] ), .S0(n3015), .S1(n3305), .Y(N246) );
  MX4XL U3003 ( .A(\IM_D_t[0][4] ), .B(\IM_D_t[1][4] ), .C(\IM_D_t[2][4] ), 
        .D(\IM_D_t[3][4] ), .S0(n3015), .S1(n3305), .Y(N247) );
  MX4XL U3004 ( .A(\IM_D_t[0][3] ), .B(\IM_D_t[1][3] ), .C(\IM_D_t[2][3] ), 
        .D(\IM_D_t[3][3] ), .S0(n3015), .S1(n3305), .Y(N248) );
  MX4XL U3005 ( .A(\IM_D_t[0][2] ), .B(\IM_D_t[1][2] ), .C(\IM_D_t[2][2] ), 
        .D(\IM_D_t[3][2] ), .S0(n3015), .S1(n3305), .Y(N249) );
  MX4XL U3006 ( .A(\IM_D_t[0][1] ), .B(\IM_D_t[1][1] ), .C(\IM_D_t[2][1] ), 
        .D(\IM_D_t[3][1] ), .S0(n3015), .S1(n3305), .Y(N250) );
  XOR2X1 U3007 ( .A(n3115), .B(n3157), .Y(N6421) );
  XNOR2XL U3008 ( .A(sec[5]), .B(n3098), .Y(N6341) );
  XNOR2XL U3009 ( .A(sec[5]), .B(\sub_819/carry[5] ), .Y(N6314) );
  XNOR2XL U3010 ( .A(sec[5]), .B(n3099), .Y(N6368) );
  XOR2XL U3011 ( .A(sec[5]), .B(\sub_825/carry[5] ), .Y(N6395) );
  XOR2X1 U3012 ( .A(n4864), .B(n3145), .Y(N6180) );
  XNOR2X1 U3013 ( .A(min[5]), .B(n3100), .Y(N6100) );
  XNOR2X1 U3014 ( .A(min[5]), .B(\sub_791/carry[5] ), .Y(N6073) );
  XNOR2X1 U3015 ( .A(min[5]), .B(n3101), .Y(N6127) );
  XOR2X1 U3016 ( .A(min[5]), .B(\sub_797/carry[5] ), .Y(N6154) );
  XOR2X1 U3017 ( .A(hour[5]), .B(n3153), .Y(N5930) );
  XNOR2X1 U3018 ( .A(hour[5]), .B(\sub_767/carry[5] ), .Y(N5904) );
  NAND2X1 U3019 ( .A(n4861), .B(n3151), .Y(\sub_767/carry[5] ) );
  NAND2X1 U3020 ( .A(n3079), .B(\r1795/carry[7] ), .Y(n3165) );
  AND2X2 U3021 ( .A(n3079), .B(n3119), .Y(n3116) );
  NAND2X1 U3022 ( .A(n3079), .B(\r1793/carry[7] ), .Y(n3164) );
  AND2X2 U3023 ( .A(n3079), .B(\r1794/carry[7] ), .Y(n3117) );
  AND2X2 U3024 ( .A(n3077), .B(\r1778/carry[6] ), .Y(n3118) );
  OR2X1 U3025 ( .A(n3077), .B(\add_772/carry[6] ), .Y(\add_772/carry[7] ) );
  AND2X2 U3026 ( .A(n3077), .B(n3120), .Y(n3119) );
  OR2X1 U3027 ( .A(n3077), .B(\r1795/carry[6] ), .Y(\r1795/carry[7] ) );
  OR2X1 U3028 ( .A(n3077), .B(n3081), .Y(\r1794/carry[7] ) );
  OR2X1 U3029 ( .A(n3077), .B(n3121), .Y(\r1793/carry[7] ) );
  OR2X1 U3030 ( .A(n3081), .B(n3075), .Y(\r1778/carry[6] ) );
  OR2X1 U3031 ( .A(n3081), .B(n3075), .Y(\add_772/carry[6] ) );
  AND2X2 U3032 ( .A(n3081), .B(\r1777/carry[5] ), .Y(n3120) );
  OR2X1 U3033 ( .A(n3081), .B(\r1795/carry[5] ), .Y(\r1795/carry[6] ) );
  AND2X2 U3034 ( .A(n3081), .B(n3122), .Y(n3121) );
  AND2X2 U3035 ( .A(n3075), .B(n3016), .Y(n3122) );
  OR2X1 U3036 ( .A(n3075), .B(n3016), .Y(\r1777/carry[5] ) );
  OR2X1 U3037 ( .A(n3075), .B(n3016), .Y(\r1795/carry[5] ) );
  XOR2X1 U3038 ( .A(n3016), .B(N6401), .Y(N6302) );
  XOR2X1 U3039 ( .A(n3016), .B(N6401), .Y(N6329) );
  XOR2X1 U3040 ( .A(n3016), .B(N6401), .Y(N6356) );
  XOR2X1 U3041 ( .A(n3016), .B(N6401), .Y(N6436) );
  XOR2X1 U3042 ( .A(n3016), .B(N6401), .Y(N6410) );
  XOR2X1 U3043 ( .A(n3016), .B(N6160), .Y(N6061) );
  XOR2X1 U3044 ( .A(n3016), .B(N6160), .Y(N6088) );
  XOR2X1 U3045 ( .A(n3016), .B(N6160), .Y(N6115) );
  XOR2X1 U3046 ( .A(n3016), .B(N6160), .Y(N6195) );
  XOR2X1 U3047 ( .A(n3016), .B(N6160), .Y(N6169) );
  XOR2X1 U3048 ( .A(n3015), .B(N1382), .Y(N1442) );
  XOR2X1 U3049 ( .A(n3015), .B(N4325), .Y(N4365) );
  XOR2X1 U3050 ( .A(n3015), .B(N7684), .Y(N4177) );
  XOR2X1 U3051 ( .A(n3015), .B(N7704), .Y(N4455) );
  XOR2X1 U3052 ( .A(n3015), .B(N670), .Y(N710) );
  XOR2X1 U3053 ( .A(n3015), .B(N2811), .Y(N2851) );
  CLKBUFX3 U3054 ( .A(n3141), .Y(n3140) );
  CLKBUFX3 U3055 ( .A(n1425), .Y(n3141) );
  XOR2X1 U3056 ( .A(N2423), .B(n2972), .Y(N3751) );
  XOR2X1 U3057 ( .A(N2422), .B(n3105), .Y(N3750) );
  XOR2X1 U3058 ( .A(N2421), .B(n3106), .Y(N3749) );
  XOR2X1 U3059 ( .A(N2420), .B(n3107), .Y(N3748) );
  XOR2X1 U3060 ( .A(N2419), .B(n3108), .Y(N3747) );
  XOR2X1 U3061 ( .A(N2418), .B(n3109), .Y(N3746) );
  XOR2X1 U3062 ( .A(N2417), .B(n3110), .Y(N3745) );
  XOR2X1 U3063 ( .A(N2416), .B(n3111), .Y(N3744) );
  XOR2X1 U3064 ( .A(N2415), .B(n3112), .Y(N3743) );
  XOR2X1 U3065 ( .A(N2414), .B(N2413), .Y(N3742) );
  CLKINVX1 U3066 ( .A(N2413), .Y(N3741) );
  XNOR2X1 U3067 ( .A(count[7]), .B(n3113), .Y(N6489) );
  XOR2X1 U3068 ( .A(count[6]), .B(n3114), .Y(N6488) );
  XOR2X1 U3069 ( .A(count[5]), .B(\add_3_root_add_0_root_add_869_4/carry[5] ), 
        .Y(N6487) );
  XNOR2X1 U3070 ( .A(count[4]), .B(count[3]), .Y(N6486) );
  MX4XL U3071 ( .A(\IM_D_t[0][23] ), .B(\IM_D_t[1][23] ), .C(\IM_D_t[2][23] ), 
        .D(\IM_D_t[3][23] ), .S0(n3015), .S1(n3305), .Y(N228) );
  MX4XL U3072 ( .A(\IM_D_t[0][22] ), .B(\IM_D_t[1][22] ), .C(\IM_D_t[2][22] ), 
        .D(\IM_D_t[3][22] ), .S0(n3015), .S1(n3305), .Y(N229) );
  MX4XL U3073 ( .A(\IM_D_t[0][21] ), .B(\IM_D_t[1][21] ), .C(\IM_D_t[2][21] ), 
        .D(\IM_D_t[3][21] ), .S0(n3015), .S1(n3305), .Y(N230) );
  MX4XL U3074 ( .A(\IM_D_t[0][20] ), .B(\IM_D_t[1][20] ), .C(\IM_D_t[2][20] ), 
        .D(\IM_D_t[3][20] ), .S0(n3015), .S1(n3305), .Y(N231) );
  MX4XL U3075 ( .A(\IM_D_t[0][19] ), .B(\IM_D_t[1][19] ), .C(\IM_D_t[2][19] ), 
        .D(\IM_D_t[3][19] ), .S0(n3015), .S1(n3305), .Y(N232) );
  MX4XL U3076 ( .A(\IM_D_t[0][18] ), .B(\IM_D_t[1][18] ), .C(\IM_D_t[2][18] ), 
        .D(\IM_D_t[3][18] ), .S0(n3015), .S1(n3305), .Y(N233) );
  MX4XL U3077 ( .A(\IM_D_t[0][17] ), .B(\IM_D_t[1][17] ), .C(\IM_D_t[2][17] ), 
        .D(\IM_D_t[3][17] ), .S0(n3015), .S1(n3305), .Y(N234) );
  MX4XL U3078 ( .A(\IM_D_t[0][16] ), .B(\IM_D_t[1][16] ), .C(\IM_D_t[2][16] ), 
        .D(\IM_D_t[3][16] ), .S0(n3015), .S1(n3305), .Y(N235) );
  MX4XL U3079 ( .A(\IM_D_t[0][15] ), .B(\IM_D_t[1][15] ), .C(\IM_D_t[2][15] ), 
        .D(\IM_D_t[3][15] ), .S0(n3015), .S1(n3305), .Y(N236) );
  MX4XL U3080 ( .A(\IM_D_t[0][14] ), .B(\IM_D_t[1][14] ), .C(\IM_D_t[2][14] ), 
        .D(\IM_D_t[3][14] ), .S0(n3015), .S1(n3305), .Y(N237) );
  MX4XL U3081 ( .A(\IM_D_t[0][13] ), .B(\IM_D_t[1][13] ), .C(\IM_D_t[2][13] ), 
        .D(\IM_D_t[3][13] ), .S0(n3015), .S1(n3305), .Y(N238) );
  MX4XL U3082 ( .A(\IM_D_t[0][12] ), .B(\IM_D_t[1][12] ), .C(\IM_D_t[2][12] ), 
        .D(\IM_D_t[3][12] ), .S0(n3015), .S1(n3305), .Y(N239) );
  MX4XL U3083 ( .A(\IM_D_t[0][11] ), .B(\IM_D_t[1][11] ), .C(\IM_D_t[2][11] ), 
        .D(\IM_D_t[3][11] ), .S0(n3015), .S1(n3305), .Y(N240) );
  MX4XL U3084 ( .A(\IM_D_t[0][10] ), .B(\IM_D_t[1][10] ), .C(\IM_D_t[2][10] ), 
        .D(\IM_D_t[3][10] ), .S0(n3015), .S1(n3305), .Y(N241) );
  MX4XL U3085 ( .A(\IM_D_t[0][9] ), .B(\IM_D_t[1][9] ), .C(\IM_D_t[2][9] ), 
        .D(\IM_D_t[3][9] ), .S0(n3015), .S1(n3305), .Y(N242) );
  XOR2X1 U3086 ( .A(n3123), .B(n3163), .Y(N5865) );
  NAND2X1 U3087 ( .A(n3079), .B(n3118), .Y(n3163) );
  XOR2X1 U3088 ( .A(n3073), .B(\add_772/carry[8] ), .Y(N5968) );
  NAND2XL U3089 ( .A(n3078), .B(n3166), .Y(\add_772/carry[8] ) );
  CLKINVX1 U3090 ( .A(\add_772/carry[7] ), .Y(n3166) );
  XOR2X1 U3091 ( .A(n3123), .B(n3165), .Y(N6028) );
  XOR2X1 U3092 ( .A(n3123), .B(n3164), .Y(N6009) );
  XOR2X1 U3093 ( .A(n3079), .B(n3118), .Y(N5864) );
  XNOR2X1 U3094 ( .A(n3079), .B(\add_772/carry[7] ), .Y(N5967) );
  XOR2X1 U3095 ( .A(n3079), .B(\r1795/carry[7] ), .Y(N6027) );
  XOR2X1 U3096 ( .A(n3079), .B(n3119), .Y(N5855) );
  XOR2X1 U3097 ( .A(n3079), .B(\r1793/carry[7] ), .Y(N6008) );
  XOR2X1 U3098 ( .A(n3079), .B(\r1794/carry[7] ), .Y(N6018) );
  XOR2X1 U3099 ( .A(n3077), .B(\r1778/carry[6] ), .Y(N5863) );
  XNOR2X1 U3100 ( .A(n3077), .B(\add_772/carry[6] ), .Y(N5966) );
  XNOR2X1 U3101 ( .A(n3077), .B(\r1795/carry[6] ), .Y(N6026) );
  XOR2X1 U3102 ( .A(n3077), .B(n3120), .Y(N5854) );
  XNOR2X1 U3103 ( .A(n3077), .B(n3121), .Y(N6007) );
  XNOR2X1 U3104 ( .A(n3077), .B(n3081), .Y(N6017) );
  XOR2X1 U3105 ( .A(n3081), .B(n3122), .Y(N6006) );
  XNOR2X1 U3106 ( .A(n3081), .B(n3075), .Y(N5965) );
  XNOR2X1 U3107 ( .A(n3081), .B(n3075), .Y(N5862) );
  XNOR2X1 U3108 ( .A(n3081), .B(\r1795/carry[5] ), .Y(N6025) );
  XOR2X1 U3109 ( .A(n3081), .B(\r1777/carry[5] ), .Y(N5853) );
  XNOR2X1 U3110 ( .A(n3075), .B(n3016), .Y(N6024) );
  XNOR2X1 U3111 ( .A(n3075), .B(n3016), .Y(N5852) );
  XOR2X1 U3112 ( .A(n3075), .B(n3016), .Y(N6005) );
  XOR2X1 U3113 ( .A(n3016), .B(N6401), .Y(N6383) );
  XOR2X1 U3114 ( .A(n3016), .B(N6160), .Y(N6142) );
  XOR2X1 U3115 ( .A(n3016), .B(N5910), .Y(N5945) );
  XOR2X1 U3116 ( .A(n3016), .B(N5910), .Y(N5919) );
  XOR2X1 U3117 ( .A(n3016), .B(N5910), .Y(N5892) );
  CLKBUFX3 U3118 ( .A(n3136), .Y(n3134) );
  CLKBUFX3 U3119 ( .A(n3139), .Y(n3137) );
  CLKBUFX3 U3120 ( .A(n3140), .Y(n3136) );
  CLKBUFX3 U3121 ( .A(n3140), .Y(n3135) );
  XOR2X1 U3122 ( .A(n3015), .B(N7622), .Y(N5022) );
  CLKBUFX3 U3123 ( .A(n3141), .Y(n3139) );
  CLKBUFX3 U3124 ( .A(n3134), .Y(n3132) );
  CLKBUFX3 U3125 ( .A(n3137), .Y(n3126) );
  CLKBUFX3 U3126 ( .A(n3138), .Y(n3133) );
  CLKBUFX3 U3127 ( .A(n3136), .Y(n3129) );
  CLKBUFX3 U3128 ( .A(n3135), .Y(n3131) );
  CLKBUFX3 U3129 ( .A(n3137), .Y(n3127) );
  CLKBUFX3 U3130 ( .A(n3136), .Y(n3128) );
  CLKBUFX3 U3131 ( .A(n3135), .Y(n3130) );
  CLKBUFX3 U3132 ( .A(n3139), .Y(n3125) );
  CLKBUFX3 U3133 ( .A(n3138), .Y(n3124) );
  CLKBUFX3 U3134 ( .A(n3139), .Y(n3138) );
  XOR2X1 U3135 ( .A(\mult_797/n2 ), .B(N6154), .Y(n3144) );
  XOR2X1 U3136 ( .A(N6153), .B(n3144), .Y(N6165) );
  XOR2X1 U3137 ( .A(\mult_799/n2 ), .B(N6180), .Y(n3146) );
  XOR2X1 U3138 ( .A(N6179), .B(n3146), .Y(N6191) );
  XOR2X1 U3139 ( .A(\mult_795/n2 ), .B(N6127), .Y(n3147) );
  XOR2X1 U3140 ( .A(N6126), .B(n3147), .Y(N6138) );
  XOR2X1 U3141 ( .A(\mult_793/n2 ), .B(N6100), .Y(n3148) );
  XOR2X1 U3142 ( .A(N6099), .B(n3148), .Y(N6111) );
  XOR2X1 U3143 ( .A(\mult_791/n2 ), .B(N6073), .Y(n3149) );
  XOR2X1 U3144 ( .A(N6072), .B(n3149), .Y(N6084) );
  XOR2X1 U3145 ( .A(\mult_789/n2 ), .B(min[5]), .Y(n3150) );
  XOR2X1 U3146 ( .A(min[4]), .B(n3150), .Y(N6057) );
  XOR2X1 U3147 ( .A(\mult_767/n2 ), .B(N5904), .Y(n3152) );
  XOR2X1 U3148 ( .A(N5903), .B(n3152), .Y(N5915) );
  XOR2X1 U3149 ( .A(\mult_769/n2 ), .B(N5930), .Y(n3154) );
  XOR2X1 U3150 ( .A(N5929), .B(n3154), .Y(N5941) );
  XOR2X1 U3151 ( .A(\mult_765/n2 ), .B(hour[5]), .Y(n3155) );
  XOR2X1 U3152 ( .A(hour[4]), .B(n3155), .Y(N5888) );
  XOR2X1 U3153 ( .A(\mult_825/n2 ), .B(N6395), .Y(n3156) );
  XOR2X1 U3154 ( .A(N6394), .B(n3156), .Y(N6406) );
  XOR2X1 U3155 ( .A(\mult_827/n2 ), .B(N6421), .Y(n3158) );
  XOR2X1 U3156 ( .A(N6420), .B(n3158), .Y(N6432) );
  XOR2X1 U3157 ( .A(\mult_823/n2 ), .B(N6368), .Y(n3159) );
  XOR2X1 U3158 ( .A(N6367), .B(n3159), .Y(N6379) );
  XOR2X1 U3159 ( .A(\mult_821/n2 ), .B(N6341), .Y(n3160) );
  XOR2X1 U3160 ( .A(N6340), .B(n3160), .Y(N6352) );
  XOR2X1 U3161 ( .A(\mult_819/n2 ), .B(N6314), .Y(n3161) );
  XOR2X1 U3162 ( .A(N6313), .B(n3161), .Y(N6325) );
  XOR2X1 U3163 ( .A(\mult_817/n2 ), .B(sec[5]), .Y(n3162) );
  XOR2X1 U3164 ( .A(sec[4]), .B(n3162), .Y(N6298) );
  OR2X1 U3165 ( .A(cycle[19]), .B(cycle[18]), .Y(n3167) );
  NOR3X1 U3166 ( .A(n3167), .B(cycle[15]), .C(cycle[14]), .Y(n3175) );
  AOI21X1 U3167 ( .A0(cycle[17]), .A1(cycle[16]), .B0(n3167), .Y(n3174) );
  NOR2X1 U3168 ( .A(cycle[13]), .B(cycle[12]), .Y(n3172) );
  NAND2X1 U3169 ( .A(cycle[11]), .B(cycle[10]), .Y(n3171) );
  OR2X1 U3170 ( .A(cycle[6]), .B(cycle[7]), .Y(n3169) );
  CLKINVX1 U3171 ( .A(n3172), .Y(n3168) );
  AOI211X1 U3172 ( .A0(cycle[8]), .A1(n3169), .B0(n3168), .C0(cycle[9]), .Y(
        n3170) );
  AOI211X1 U3173 ( .A0(n3172), .A1(n3171), .B0(n3170), .C0(n3174), .Y(n3173)
         );
  AOI2BB1X1 U3174 ( .A0N(n3177), .A1N(n3176), .B0(offset_w[15]), .Y(N2136) );
  NAND4X1 U3175 ( .A(N798), .B(n3073), .C(N800), .D(N799), .Y(n3179) );
  NAND2X1 U3176 ( .A(N802), .B(N801), .Y(n3178) );
  AO22X1 U3177 ( .A0(n3180), .A1(n3179), .B0(n3180), .B1(n3178), .Y(N3841) );
  XOR2X1 U3178 ( .A(tick[0]), .B(n3181), .Y(n1689) );
  CLKMX2X2 U3179 ( .A(n3182), .B(n3183), .S0(n2980), .Y(n1688) );
  MXI2X1 U3180 ( .A(n3184), .B(n3185), .S0(tick[2]), .Y(n1687) );
  NOR2X1 U3181 ( .A(n2980), .B(n3182), .Y(n3185) );
  OAI21XL U3182 ( .A0(tick[0]), .A1(n3186), .B0(n3181), .Y(n3182) );
  NAND2X1 U3183 ( .A(n3183), .B(tick[1]), .Y(n3184) );
  NOR2BX1 U3184 ( .AN(tick[0]), .B(n3187), .Y(n3183) );
  AO22X1 U3185 ( .A0(n3188), .A1(n3189), .B0(n144), .B1(n3190), .Y(n1686) );
  NAND4BX1 U3186 ( .AN(n3191), .B(n3192), .C(n3193), .D(n3194), .Y(n1685) );
  AOI221XL U3187 ( .A0(n3195), .A1(N3732), .B0(n3196), .B1(IM_A[0]), .C0(n3198), .Y(n3194) );
  OAI21XL U3188 ( .A0(n1424), .A1(n3199), .B0(n3200), .Y(n3198) );
  NOR2X1 U3189 ( .A(n3205), .B(n3206), .Y(n3204) );
  CLKINVX1 U3190 ( .A(n3207), .Y(n3203) );
  AOI222XL U3191 ( .A0(n3208), .A1(n3209), .B0(n3210), .B1(n3211), .C0(n3212), 
        .C1(n3213), .Y(n3193) );
  NAND4X1 U3192 ( .A(n3214), .B(n3215), .C(n3216), .D(n3217), .Y(n3213) );
  AOI222XL U3193 ( .A0(N3752), .A1(n3218), .B0(n3219), .B1(IM_A[0]), .C0(N3617), .C1(n3220), .Y(n3217) );
  AOI22X1 U3194 ( .A0(N3732), .A1(n3221), .B0(N3732), .B1(n3222), .Y(n3216) );
  NAND4X1 U3195 ( .A(n3227), .B(n3228), .C(n3229), .D(n3230), .Y(n3211) );
  AOI222XL U3196 ( .A0(n3231), .A1(N1024), .B0(N867), .B1(n3232), .C0(n3233), 
        .C1(IM_A[0]), .Y(n3230) );
  AOI22X1 U3197 ( .A0(N807), .A1(n3234), .B0(N1279), .B1(n3235), .Y(n3229) );
  AOI22X1 U3198 ( .A0(n3236), .A1(N487), .B0(N1356), .B1(n3237), .Y(n3228) );
  AOI222XL U3199 ( .A0(N6550), .A1(n3240), .B0(n3241), .B1(n3242), .C0(n3243), 
        .C1(N2318), .Y(n3192) );
  OAI222XL U3200 ( .A0(n3244), .A1(n3245), .B0(n3246), .B1(n3247), .C0(n3248), 
        .C1(n3249), .Y(n3191) );
  AND4X1 U3201 ( .A(n3250), .B(n3251), .C(n3252), .D(n3253), .Y(n3245) );
  AOI222XL U3202 ( .A0(N508), .A1(n3254), .B0(N487), .B1(n3255), .C0(n3256), 
        .C1(IM_A[0]), .Y(n3253) );
  AOI22X1 U3203 ( .A0(N548), .A1(n3257), .B0(n3232), .B1(N1024), .Y(n3252) );
  CLKINVX1 U3204 ( .A(n3258), .Y(n3232) );
  AOI222XL U3205 ( .A0(N644), .A1(n3237), .B0(N867), .B1(n3231), .C0(N944), 
        .C1(n3234), .Y(n3251) );
  CLKINVX1 U3206 ( .A(n3259), .Y(n3231) );
  AOI22X1 U3207 ( .A0(N709), .A1(n3238), .B0(N807), .B1(n3239), .Y(n3250) );
  AO22X1 U3208 ( .A0(N6483), .A1(n3189), .B0(n143), .B1(n3190), .Y(n1684) );
  NOR4X1 U3209 ( .A(n3264), .B(n3265), .C(n3266), .D(n3267), .Y(n3263) );
  AO22X1 U3210 ( .A0(n3212), .A1(n3268), .B0(n3210), .B1(n3269), .Y(n3267) );
  AOI222XL U3211 ( .A0(N1357), .A1(n3237), .B0(N1280), .B1(n3235), .C0(N488), 
        .C1(n3236), .Y(n3273) );
  NAND4X1 U3212 ( .A(n3274), .B(n3275), .C(n3276), .D(n3277), .Y(n3268) );
  AOI222XL U3213 ( .A0(N3753), .A1(n3218), .B0(n3219), .B1(IM_A[1]), .C0(N3618), .C1(n3220), .Y(n3277) );
  AOI22X1 U3214 ( .A0(N3733), .A1(n3221), .B0(N3733), .B1(n3222), .Y(n3276) );
  OAI22XL U3215 ( .A0(n3279), .A1(n3244), .B0(n3280), .B1(n3248), .Y(n3266) );
  AOI211X1 U3216 ( .A0(N645), .A1(n3237), .B0(n3281), .C0(n3282), .Y(n3279) );
  AO22X1 U3217 ( .A0(N549), .A1(n3257), .B0(N509), .B1(n3254), .Y(n3282) );
  OAI2BB2XL U3218 ( .B0(n3283), .B1(n3246), .A0N(N3733), .A1N(n3195), .Y(n3265) );
  OAI222XL U3219 ( .A0(n3284), .A1(n3285), .B0(n4875), .B1(n3199), .C0(n3286), 
        .C1(n3271), .Y(n3264) );
  CLKINVX1 U3220 ( .A(N945), .Y(n3271) );
  CLKINVX1 U3221 ( .A(N808), .Y(n3285) );
  AOI211X1 U3222 ( .A0(N6551), .A1(n3240), .B0(n3287), .C0(n3288), .Y(n3262)
         );
  MXI2X1 U3223 ( .A(n3200), .B(n3289), .S0(n4788), .Y(n3288) );
  OAI2BB2XL U3224 ( .B0(n4843), .B1(n3290), .A0N(N2319), .A1N(n3243), .Y(n3287) );
  AOI22X1 U3225 ( .A0(N868), .A1(n3291), .B0(N1025), .B1(n3292), .Y(n3261) );
  OAI222XL U3226 ( .A0(n3293), .A1(n3294), .B0(n3295), .B1(n3296), .C0(n3297), 
        .C1(n3298), .Y(n3260) );
  CLKINVX1 U3227 ( .A(N488), .Y(n3294) );
  AO22X1 U3228 ( .A0(N6484), .A1(n3189), .B0(n142), .B1(n3190), .Y(n1682) );
  MXI2X1 U3229 ( .A(n2965), .B(n3299), .S0(n3300), .Y(n1681) );
  MXI2X1 U3230 ( .A(n3301), .B(n3302), .S0(n4854), .Y(n1680) );
  MXI2X1 U3231 ( .A(n3303), .B(n3304), .S0(n4856), .Y(n1679) );
  NAND3X1 U3232 ( .A(n3305), .B(n3306), .C(n3307), .Y(n3304) );
  MXI2X1 U3233 ( .A(n3308), .B(n3309), .S0(n4855), .Y(n1678) );
  NAND2X1 U3234 ( .A(n3307), .B(n3306), .Y(n3309) );
  OAI21XL U3235 ( .A0(n3310), .A1(n4743), .B0(n3311), .Y(n1677) );
  AOI22X1 U3236 ( .A0(N4631), .A1(n3312), .B0(n86), .B1(n3313), .Y(n3311) );
  OAI21XL U3237 ( .A0(n3310), .A1(n4737), .B0(n3314), .Y(n1676) );
  AOI22X1 U3238 ( .A0(N4646), .A1(n3312), .B0(n71), .B1(n3313), .Y(n3314) );
  OAI211X1 U3239 ( .A0(n3315), .A1(n3316), .B0(n3317), .C0(n3318), .Y(n1675)
         );
  AOI222XL U3240 ( .A0(n3319), .A1(n3320), .B0(n3321), .B1(n3322), .C0(n3323), 
        .C1(n3324), .Y(n3318) );
  NOR2X1 U3241 ( .A(n3186), .B(n3325), .Y(n3323) );
  OAI221XL U3242 ( .A0(n3326), .A1(n3327), .B0(n3328), .B1(n3329), .C0(n3330), 
        .Y(n3320) );
  NAND3BX1 U3243 ( .AN(n3331), .B(n3332), .C(n3333), .Y(n3330) );
  NAND3X1 U3244 ( .A(n3334), .B(n3335), .C(n3336), .Y(n3327) );
  NAND3X1 U3245 ( .A(n3337), .B(n3338), .C(n3339), .Y(n3326) );
  OAI21XL U3246 ( .A0(n3340), .A1(n3341), .B0(state[2]), .Y(n3317) );
  AOI221XL U3247 ( .A0(n3342), .A1(n3343), .B0(n3344), .B1(n3345), .C0(n3346), 
        .Y(n3315) );
  NOR3X1 U3248 ( .A(n3347), .B(N3841), .C(n3348), .Y(n3346) );
  CLKINVX1 U3249 ( .A(n3349), .Y(n3345) );
  NAND3X1 U3250 ( .A(n3350), .B(n3351), .C(n3352), .Y(n1674) );
  AOI222XL U3251 ( .A0(n3353), .A1(n3354), .B0(state[0]), .B1(n3355), .C0(
        n3356), .C1(n3357), .Y(n3352) );
  CLKINVX1 U3252 ( .A(n3358), .Y(n3355) );
  AOI211X1 U3253 ( .A0(n3359), .A1(n3360), .B0(n3361), .C0(n3341), .Y(n3358)
         );
  OAI221XL U3254 ( .A0(n3362), .A1(n3363), .B0(n3364), .B1(n3365), .C0(n3366), 
        .Y(n3341) );
  AOI211X1 U3255 ( .A0(n3367), .A1(n3368), .B0(n3369), .C0(n3357), .Y(n3366)
         );
  NAND3X1 U3256 ( .A(n3324), .B(n3370), .C(n3186), .Y(n3351) );
  AOI32X1 U3257 ( .A0(n3371), .A1(n3372), .A2(n2964), .B0(n3373), .B1(n3374), 
        .Y(n3350) );
  OAI222XL U3258 ( .A0(n3375), .A1(n3376), .B0(n3377), .B1(n3378), .C0(n3379), 
        .C1(n3244), .Y(n3374) );
  AO22X1 U3259 ( .A0(n3380), .A1(n3381), .B0(n3332), .B1(n3382), .Y(n1673) );
  OAI32X1 U3260 ( .A0(n3328), .A1(n3202), .A2(n3381), .B0(n3316), .B1(n3383), 
        .Y(n3382) );
  OAI211X1 U3261 ( .A0(n3384), .A1(n3385), .B0(n3386), .C0(n3387), .Y(n3380)
         );
  AOI211X1 U3262 ( .A0(n3388), .A1(n3389), .B0(n3390), .C0(n3391), .Y(n3387)
         );
  NAND2X1 U3263 ( .A(n3362), .B(n3392), .Y(n3389) );
  NOR4BX1 U3264 ( .AN(n3393), .B(n4706), .C(n4705), .D(n3394), .Y(n3362) );
  NOR4X1 U3265 ( .A(n4701), .B(n4702), .C(n4703), .D(n4704), .Y(n3393) );
  OAI21XL U3266 ( .A0(n3186), .A1(n3325), .B0(n3363), .Y(n3388) );
  NOR2X1 U3267 ( .A(n3395), .B(n3396), .Y(n3385) );
  OAI21XL U3268 ( .A0(n3310), .A1(n4736), .B0(n3397), .Y(n1672) );
  AOI22X1 U3269 ( .A0(N4632), .A1(n3312), .B0(n85), .B1(n3313), .Y(n3397) );
  OAI21XL U3270 ( .A0(n3310), .A1(n4738), .B0(n3398), .Y(n1671) );
  AOI22X1 U3271 ( .A0(N4645), .A1(n3312), .B0(n72), .B1(n3313), .Y(n3398) );
  NAND4X1 U3272 ( .A(n3378), .B(n3399), .C(n3400), .D(n3401), .Y(n1670) );
  AOI211X1 U3273 ( .A0(n3367), .A1(n3368), .B0(n3402), .C0(n3403), .Y(n3401)
         );
  OA21XL U3274 ( .A0(N3841), .A1(n3348), .B0(n3372), .Y(n3404) );
  NAND3X1 U3275 ( .A(n3406), .B(n3407), .C(n3363), .Y(n3402) );
  CLKINVX1 U3276 ( .A(n3321), .Y(n3363) );
  NOR2X1 U3277 ( .A(n3325), .B(n3324), .Y(n3321) );
  NAND2X1 U3278 ( .A(n3201), .B(n3408), .Y(n3368) );
  AOI221XL U3279 ( .A0(n3319), .A1(n3409), .B0(n3410), .B1(n3411), .C0(n3412), 
        .Y(n3400) );
  NOR3BXL U3280 ( .AN(n3413), .B(n3348), .C(n3414), .Y(n3412) );
  OAI22XL U3281 ( .A0(n3342), .A1(n3415), .B0(n3344), .B1(n3349), .Y(n3411) );
  OAI211X1 U3282 ( .A0(n3416), .A1(n3417), .B0(n3418), .C0(n3419), .Y(n3409)
         );
  CLKINVX1 U3283 ( .A(n3420), .Y(n3419) );
  OAI21XL U3284 ( .A0(N2136), .A1(n3421), .B0(n3422), .Y(n3418) );
  NAND2X1 U3285 ( .A(n3364), .B(n3423), .Y(n3399) );
  NOR2X1 U3286 ( .A(n3210), .B(n3371), .Y(n3378) );
  AO22X1 U3287 ( .A0(count[3]), .A1(n3189), .B0(n141), .B1(n3190), .Y(n1669)
         );
  AO22X1 U3288 ( .A0(count[4]), .A1(n3189), .B0(n140), .B1(n3190), .Y(n1668)
         );
  AO22X1 U3289 ( .A0(n3424), .A1(n3189), .B0(n139), .B1(n3190), .Y(n1667) );
  AO22X1 U3290 ( .A0(n3425), .A1(n3189), .B0(n138), .B1(n3190), .Y(n1666) );
  AO22X1 U3291 ( .A0(n3426), .A1(n3189), .B0(n137), .B1(n3190), .Y(n1665) );
  OAI31XL U3292 ( .A0(n3428), .A1(n3429), .A2(n3430), .B0(n3431), .Y(n3427) );
  OAI2BB2XL U3293 ( .B0(n3364), .B1(n3365), .A0N(n3432), .A1N(n3433), .Y(n3430) );
  OAI22XL U3294 ( .A0(n3316), .A1(n3434), .B0(n3435), .B1(n3436), .Y(n3429) );
  CLKINVX1 U3295 ( .A(n3437), .Y(n3428) );
  AOI211X1 U3296 ( .A0(n3438), .A1(n3357), .B0(n3361), .C0(n3439), .Y(n3437)
         );
  OAI32X1 U3297 ( .A0(n3440), .A1(n3441), .A2(n3442), .B0(n3199), .B1(n3353), 
        .Y(n3439) );
  AOI21X1 U3298 ( .A0(n3445), .A1(n3319), .B0(n3446), .Y(n3444) );
  AOI31X1 U3299 ( .A0(n3447), .A1(n3448), .A2(n3449), .B0(n3359), .Y(n3443) );
  OAI21XL U3300 ( .A0(n3450), .A1(n3451), .B0(n3452), .Y(n3359) );
  OAI22XL U3301 ( .A0(n3302), .A1(n3348), .B0(n4857), .B1(n3453), .Y(n1664) );
  OA21XL U3302 ( .A0(n3302), .A1(\gt_332/n15 ), .B0(n3303), .Y(n3453) );
  OA21XL U3303 ( .A0(n3302), .A1(n3305), .B0(n3308), .Y(n3303) );
  OA21XL U3304 ( .A0(n3302), .A1(n3306), .B0(n3301), .Y(n3308) );
  NOR4X1 U3305 ( .A(n3361), .B(n3390), .C(n3454), .D(n3455), .Y(n3301) );
  OAI221XL U3306 ( .A0(n3456), .A1(n3457), .B0(n3201), .B1(n3458), .C0(n3459), 
        .Y(n3455) );
  OAI21XL U3307 ( .A0(n3384), .A1(n3415), .B0(n3460), .Y(n3454) );
  CLKINVX1 U3308 ( .A(n3461), .Y(n3361) );
  CLKINVX1 U3309 ( .A(n3307), .Y(n3302) );
  AOI32X1 U3310 ( .A0(n3456), .A1(n3348), .A2(n3413), .B0(n3445), .B1(n3465), 
        .Y(n3464) );
  NAND2X1 U3311 ( .A(n3440), .B(n3316), .Y(n3465) );
  CLKINVX1 U3312 ( .A(n3414), .Y(n3456) );
  NOR2X1 U3313 ( .A(n3468), .B(n3469), .Y(n3377) );
  CLKMX2X2 U3314 ( .A(pic_size[6]), .B(IM_Q[6]), .S0(n3300), .Y(n1661) );
  CLKMX2X2 U3315 ( .A(pic_size[5]), .B(IM_Q[5]), .S0(n3300), .Y(n1660) );
  CLKMX2X2 U3316 ( .A(pic_size[4]), .B(IM_Q[4]), .S0(n3300), .Y(n1659) );
  CLKMX2X2 U3317 ( .A(pic_size[3]), .B(IM_Q[3]), .S0(n3300), .Y(n1658) );
  OAI31XL U3318 ( .A0(n3477), .A1(n3478), .A2(n3479), .B0(n3480), .Y(n1654) );
  OAI31XL U3319 ( .A0(n3481), .A1(n3478), .A2(n3482), .B0(n2979), .Y(n3480) );
  NAND3X1 U3320 ( .A(n3483), .B(n3415), .C(n3332), .Y(n3481) );
  OAI211X1 U3321 ( .A0(n3484), .A1(n3082), .B0(n3485), .C0(n3486), .Y(n1653)
         );
  AOI222XL U3322 ( .A0(N2944), .A1(n3487), .B0(N2488), .B1(n3488), .C0(N4615), 
        .C1(n3489), .Y(n3486) );
  AOI22X1 U3323 ( .A0(N3213), .A1(n3490), .B0(n102), .B1(n3491), .Y(n3485) );
  AOI222XL U3324 ( .A0(N2954), .A1(n3487), .B0(N2498), .B1(n3488), .C0(N4625), 
        .C1(n3489), .Y(n3493) );
  AOI222XL U3325 ( .A0(N2959), .A1(n3487), .B0(N2503), .B1(n3488), .C0(N4630), 
        .C1(n3489), .Y(n3495) );
  AOI22X1 U3326 ( .A0(N3228), .A1(n3490), .B0(n87), .B1(n3491), .Y(n3494) );
  OAI211X1 U3327 ( .A0(n3484), .A1(n2985), .B0(n3496), .C0(n3497), .Y(n1650)
         );
  AOI222XL U3328 ( .A0(N2958), .A1(n3487), .B0(N2502), .B1(n3488), .C0(N4629), 
        .C1(n3489), .Y(n3497) );
  AOI22X1 U3329 ( .A0(N3227), .A1(n3490), .B0(n88), .B1(n3491), .Y(n3496) );
  AOI222XL U3330 ( .A0(N2957), .A1(n3487), .B0(N2501), .B1(n3488), .C0(N4628), 
        .C1(n3489), .Y(n3499) );
  AOI222XL U3331 ( .A0(N2956), .A1(n3487), .B0(N2500), .B1(n3488), .C0(N4627), 
        .C1(n3489), .Y(n3501) );
  AOI222XL U3332 ( .A0(N2955), .A1(n3487), .B0(N2499), .B1(n3488), .C0(N4626), 
        .C1(n3489), .Y(n3503) );
  AOI222XL U3333 ( .A0(N2953), .A1(n3487), .B0(N2497), .B1(n3488), .C0(N4624), 
        .C1(n3489), .Y(n3505) );
  OAI211X1 U3334 ( .A0(n3484), .A1(n3123), .B0(n3506), .C0(n3507), .Y(n1645)
         );
  AOI222XL U3335 ( .A0(N2952), .A1(n3487), .B0(N2496), .B1(n3488), .C0(N4623), 
        .C1(n3489), .Y(n3507) );
  AOI22X1 U3336 ( .A0(N3221), .A1(n3490), .B0(n94), .B1(n3491), .Y(n3506) );
  OAI211X1 U3337 ( .A0(n3484), .A1(n3078), .B0(n3508), .C0(n3509), .Y(n1644)
         );
  AOI222XL U3338 ( .A0(N2951), .A1(n3487), .B0(N2495), .B1(n3488), .C0(N4622), 
        .C1(n3489), .Y(n3509) );
  AOI22X1 U3339 ( .A0(N3220), .A1(n3490), .B0(n95), .B1(n3491), .Y(n3508) );
  OAI211X1 U3340 ( .A0(n3484), .A1(n3076), .B0(n3510), .C0(n3511), .Y(n1643)
         );
  AOI222XL U3341 ( .A0(N2950), .A1(n3487), .B0(N2494), .B1(n3488), .C0(N4621), 
        .C1(n3489), .Y(n3511) );
  AOI22X1 U3342 ( .A0(N3219), .A1(n3490), .B0(n96), .B1(n3491), .Y(n3510) );
  OAI211X1 U3343 ( .A0(n3484), .A1(n3080), .B0(n3512), .C0(n3513), .Y(n1642)
         );
  AOI222XL U3344 ( .A0(N2949), .A1(n3487), .B0(N2493), .B1(n3488), .C0(N4620), 
        .C1(n3489), .Y(n3513) );
  AOI22X1 U3345 ( .A0(N3218), .A1(n3490), .B0(n97), .B1(n3491), .Y(n3512) );
  OAI211X1 U3346 ( .A0(n3484), .A1(n3074), .B0(n3514), .C0(n3515), .Y(n1641)
         );
  AOI222XL U3347 ( .A0(N2948), .A1(n3487), .B0(N2492), .B1(n3488), .C0(N4619), 
        .C1(n3489), .Y(n3515) );
  AOI22X1 U3348 ( .A0(N3217), .A1(n3490), .B0(n98), .B1(n3491), .Y(n3514) );
  OAI211X1 U3349 ( .A0(n3484), .A1(n2982), .B0(n3516), .C0(n3517), .Y(n1640)
         );
  AOI222XL U3350 ( .A0(N2947), .A1(n3487), .B0(N2491), .B1(n3488), .C0(N4618), 
        .C1(n3489), .Y(n3517) );
  AOI22X1 U3351 ( .A0(N3216), .A1(n3490), .B0(n99), .B1(n3491), .Y(n3516) );
  OAI211X1 U3352 ( .A0(n3484), .A1(n2968), .B0(n3518), .C0(n3519), .Y(n1639)
         );
  AOI222XL U3353 ( .A0(N2946), .A1(n3487), .B0(N2490), .B1(n3488), .C0(N4617), 
        .C1(n3489), .Y(n3519) );
  AOI22X1 U3354 ( .A0(N3215), .A1(n3490), .B0(n100), .B1(n3491), .Y(n3518) );
  OAI211X1 U3355 ( .A0(n3484), .A1(n2961), .B0(n3520), .C0(n3521), .Y(n1638)
         );
  AOI222XL U3356 ( .A0(N2945), .A1(n3487), .B0(N2489), .B1(n3488), .C0(N4616), 
        .C1(n3489), .Y(n3521) );
  NOR4X1 U3357 ( .A(n3344), .B(n3527), .C(n3528), .D(n3417), .Y(n3525) );
  AOI32X1 U3358 ( .A0(n3531), .A1(n3532), .A2(n3360), .B0(n3413), .B1(n3414), 
        .Y(n3530) );
  NAND4X1 U3359 ( .A(n3533), .B(n3534), .C(n3535), .D(n3536), .Y(n3414) );
  NOR4X1 U3360 ( .A(N798), .B(n3073), .C(n3079), .D(n3077), .Y(n3536) );
  NOR4X1 U3361 ( .A(n3081), .B(n3016), .C(N804), .D(N803), .Y(n3535) );
  NOR4X1 U3362 ( .A(N802), .B(N801), .C(N800), .D(N799), .Y(n3534) );
  NOR4X1 U3363 ( .A(n3082), .B(n2961), .C(n2968), .D(n3074), .Y(n3533) );
  OAI31XL U3364 ( .A0(n3349), .A1(n3344), .A2(n3537), .B0(n3434), .Y(n3532) );
  NAND2X1 U3365 ( .A(n3395), .B(n3538), .Y(n3434) );
  CLKINVX1 U3366 ( .A(n3539), .Y(n3395) );
  CLKINVX1 U3367 ( .A(n3447), .Y(n3537) );
  CLKINVX1 U3368 ( .A(n3448), .Y(n3344) );
  NAND4X1 U3369 ( .A(n3540), .B(n3541), .C(n3542), .D(n3543), .Y(n3448) );
  NOR4X1 U3370 ( .A(n3544), .B(n3545), .C(n3546), .D(n3547), .Y(n3543) );
  XOR2X1 U3371 ( .A(N5164), .B(n3548), .Y(n3547) );
  XOR2X1 U3372 ( .A(N5166), .B(n3549), .Y(n3546) );
  XOR2X1 U3373 ( .A(N5165), .B(n3550), .Y(n3545) );
  NAND3X1 U3374 ( .A(n3551), .B(n3552), .C(n3553), .Y(n3544) );
  XOR2X1 U3375 ( .A(N5152), .B(n3554), .Y(n3553) );
  XOR2X1 U3376 ( .A(N5163), .B(n3555), .Y(n3551) );
  NOR4X1 U3377 ( .A(n3556), .B(n3557), .C(n3558), .D(n3559), .Y(n3542) );
  XNOR2X1 U3378 ( .A(N5148), .B(n3296), .Y(n3559) );
  AOI221XL U3379 ( .A0(N4977), .A1(n3560), .B0(N5022), .B1(n3561), .C0(n3562), 
        .Y(n3296) );
  XOR2X1 U3380 ( .A(N5151), .B(n3563), .Y(n3558) );
  XOR2X1 U3381 ( .A(N5147), .B(n3209), .Y(n3557) );
  CLKINVX1 U3382 ( .A(n3564), .Y(n3209) );
  AOI221XL U3383 ( .A0(N4976), .A1(n3560), .B0(N5021), .B1(n3561), .C0(n3565), 
        .Y(n3564) );
  NAND2X1 U3384 ( .A(n3566), .B(n3567), .Y(n3556) );
  XOR2X1 U3385 ( .A(N5153), .B(n3568), .Y(n3567) );
  XOR2X1 U3386 ( .A(N5154), .B(n3569), .Y(n3566) );
  NOR4X1 U3387 ( .A(n3570), .B(n3571), .C(n3572), .D(n3573), .Y(n3541) );
  XNOR2X1 U3388 ( .A(N5150), .B(n3574), .Y(n3573) );
  XOR2X1 U3389 ( .A(N5160), .B(n3575), .Y(n3572) );
  XOR2X1 U3390 ( .A(N5159), .B(n3576), .Y(n3571) );
  NAND2X1 U3391 ( .A(n3577), .B(n3578), .Y(n3570) );
  XOR2X1 U3392 ( .A(N5162), .B(n3579), .Y(n3578) );
  XOR2X1 U3393 ( .A(N5149), .B(n3580), .Y(n3577) );
  NOR4X1 U3394 ( .A(n3581), .B(n3582), .C(n3583), .D(n3584), .Y(n3540) );
  XOR2X1 U3395 ( .A(N5155), .B(n3585), .Y(n3584) );
  XOR2X1 U3396 ( .A(N5157), .B(n3586), .Y(n3583) );
  XOR2X1 U3397 ( .A(N5156), .B(n3587), .Y(n3582) );
  NAND2X1 U3398 ( .A(n3588), .B(n3589), .Y(n3581) );
  XOR2X1 U3399 ( .A(N5158), .B(n3590), .Y(n3589) );
  XOR2X1 U3400 ( .A(N5161), .B(n3591), .Y(n3588) );
  OAI21XL U3401 ( .A0(n3255), .A1(n3432), .B0(n3433), .Y(n3529) );
  OAI211X1 U3402 ( .A0(n3592), .A1(n3539), .B0(n3593), .C0(n3594), .Y(n3432)
         );
  NAND3BX1 U3403 ( .AN(n3416), .B(n3447), .C(n3449), .Y(n3594) );
  NAND4X1 U3404 ( .A(n3595), .B(n4870), .C(n4871), .D(n3188), .Y(n3447) );
  NAND2X1 U3405 ( .A(n3338), .B(n3596), .Y(n3416) );
  NAND4X1 U3406 ( .A(n3334), .B(n3335), .C(n3339), .D(n3337), .Y(n3596) );
  AND4X1 U3407 ( .A(n3597), .B(n3598), .C(n3599), .D(n3600), .Y(n3337) );
  XOR2X1 U3408 ( .A(N2993), .B(n3601), .Y(n3600) );
  NOR2X1 U3409 ( .A(n3602), .B(n3603), .Y(n3599) );
  XNOR2X1 U3410 ( .A(N2992), .B(n3604), .Y(n3603) );
  XNOR2X1 U3411 ( .A(N2994), .B(n3605), .Y(n3602) );
  XOR2X1 U3412 ( .A(N2995), .B(n3606), .Y(n3598) );
  XOR2X1 U3413 ( .A(N2998), .B(n3607), .Y(n3597) );
  AND4X1 U3414 ( .A(n3608), .B(n3609), .C(n3610), .D(n3611), .Y(n3339) );
  XOR2X1 U3415 ( .A(N2996), .B(n3612), .Y(n3611) );
  NOR2X1 U3416 ( .A(n3613), .B(n3614), .Y(n3610) );
  XNOR2X1 U3417 ( .A(N2987), .B(n3615), .Y(n3614) );
  XNOR2X1 U3418 ( .A(N2997), .B(n3616), .Y(n3613) );
  XOR2X1 U3419 ( .A(N2999), .B(n3617), .Y(n3609) );
  XOR2X1 U3420 ( .A(N2986), .B(n3618), .Y(n3608) );
  AND4X1 U3421 ( .A(n3619), .B(n3620), .C(n3621), .D(n3622), .Y(n3335) );
  XOR2X1 U3422 ( .A(N2984), .B(n3247), .Y(n3622) );
  AOI221XL U3423 ( .A0(N2785), .A1(n3560), .B0(N2850), .B1(n3561), .C0(n3565), 
        .Y(n3247) );
  NOR2X1 U3424 ( .A(n3623), .B(n1423), .Y(n3565) );
  NOR2X1 U3425 ( .A(n3624), .B(n3625), .Y(n3621) );
  XNOR2X1 U3426 ( .A(N2985), .B(n3283), .Y(n3625) );
  AOI221XL U3427 ( .A0(N2786), .A1(n3560), .B0(N2851), .B1(n3561), .C0(n3562), 
        .Y(n3283) );
  NOR2X1 U3428 ( .A(n3623), .B(n4843), .Y(n3562) );
  XNOR2X1 U3429 ( .A(N2988), .B(n3626), .Y(n3624) );
  XOR2X1 U3430 ( .A(N2990), .B(n3627), .Y(n3620) );
  XOR2X1 U3431 ( .A(N2991), .B(n3628), .Y(n3619) );
  AND4X1 U3432 ( .A(n3629), .B(n3630), .C(n3631), .D(n3632), .Y(n3334) );
  NOR3X1 U3433 ( .A(n3633), .B(N3004), .C(n3634), .Y(n3632) );
  XNOR2X1 U3434 ( .A(N3000), .B(n3635), .Y(n3634) );
  XNOR2X1 U3435 ( .A(N2989), .B(n3636), .Y(n3633) );
  XOR2X1 U3436 ( .A(N3002), .B(n3637), .Y(n3631) );
  XOR2X1 U3437 ( .A(N3003), .B(n3638), .Y(n3630) );
  XOR2X1 U3438 ( .A(N3001), .B(n3639), .Y(n3629) );
  OAI2BB1X1 U3439 ( .A0N(n3524), .A1N(n3483), .B0(n3421), .Y(n3593) );
  NAND2X1 U3440 ( .A(n3343), .B(n3421), .Y(n3539) );
  CLKINVX1 U3441 ( .A(n3640), .Y(n3435) );
  CLKINVX1 U3442 ( .A(n3332), .Y(n3421) );
  AOI2BB1X1 U3443 ( .A0N(n3384), .A1N(n3531), .B0(n3645), .Y(n3644) );
  OR2X1 U3444 ( .A(n3523), .B(n3450), .Y(n3643) );
  NAND2X1 U3445 ( .A(n3422), .B(n3360), .Y(n3523) );
  AO21X1 U3446 ( .A0(n3440), .A1(n3527), .B0(n3452), .Y(n3642) );
  NOR2X1 U3447 ( .A(n3445), .B(n3646), .Y(n3452) );
  CLKINVX1 U3448 ( .A(n3408), .Y(n3445) );
  NAND2X1 U3449 ( .A(n3340), .B(n3647), .Y(n3461) );
  OAI21XL U3450 ( .A0(n3310), .A1(n4739), .B0(n3648), .Y(n1637) );
  AOI22X1 U3451 ( .A0(N4644), .A1(n3312), .B0(n73), .B1(n3313), .Y(n3648) );
  OAI21XL U3452 ( .A0(n3310), .A1(n4740), .B0(n3649), .Y(n1636) );
  AOI22X1 U3453 ( .A0(N4643), .A1(n3312), .B0(n74), .B1(n3313), .Y(n3649) );
  OAI21XL U3454 ( .A0(n3310), .A1(n4741), .B0(n3650), .Y(n1635) );
  AOI22X1 U3455 ( .A0(N4642), .A1(n3312), .B0(n75), .B1(n3313), .Y(n3650) );
  OAI21XL U3456 ( .A0(n3310), .A1(n4742), .B0(n3651), .Y(n1634) );
  AOI22X1 U3457 ( .A0(N4641), .A1(n3312), .B0(n76), .B1(n3313), .Y(n3651) );
  OAI21XL U3458 ( .A0(n3310), .A1(n4728), .B0(n3652), .Y(n1633) );
  AOI22X1 U3459 ( .A0(N4640), .A1(n3312), .B0(n77), .B1(n3313), .Y(n3652) );
  OAI21XL U3460 ( .A0(n3310), .A1(n4729), .B0(n3653), .Y(n1632) );
  AOI22X1 U3461 ( .A0(N4639), .A1(n3312), .B0(n78), .B1(n3313), .Y(n3653) );
  OAI21XL U3462 ( .A0(n3310), .A1(n4730), .B0(n3654), .Y(n1631) );
  OAI21XL U3463 ( .A0(n3310), .A1(n4731), .B0(n3655), .Y(n1630) );
  OAI21XL U3464 ( .A0(n3310), .A1(n4732), .B0(n3656), .Y(n1629) );
  OAI21XL U3465 ( .A0(n3310), .A1(n4733), .B0(n3657), .Y(n1628) );
  OAI21XL U3466 ( .A0(n3310), .A1(n4734), .B0(n3658), .Y(n1627) );
  OAI21XL U3467 ( .A0(n3310), .A1(n4735), .B0(n3659), .Y(n1626) );
  CLKINVX1 U3468 ( .A(n3661), .Y(n3479) );
  MXI2X1 U3469 ( .A(n3662), .B(n3663), .S0(N444), .Y(n3660) );
  AOI21X1 U3470 ( .A0(n3531), .A1(n3664), .B0(n3420), .Y(n3663) );
  OAI21XL U3471 ( .A0(n3592), .A1(n3328), .B0(n3665), .Y(n3420) );
  CLKINVX1 U3472 ( .A(n3329), .Y(n3592) );
  NAND4X1 U3473 ( .A(n3666), .B(n3667), .C(n3668), .D(n3669), .Y(n3329) );
  NOR4X1 U3474 ( .A(n3670), .B(n3671), .C(n3672), .D(n3673), .Y(n3669) );
  XNOR2X1 U3475 ( .A(N3001), .B(n3674), .Y(n3673) );
  XNOR2X1 U3476 ( .A(N3003), .B(n3675), .Y(n3672) );
  XNOR2X1 U3477 ( .A(N3002), .B(n3676), .Y(n3671) );
  NAND3BX1 U3478 ( .AN(N3004), .B(n3677), .C(n3678), .Y(n3670) );
  XOR2X1 U3479 ( .A(n3679), .B(N2989), .Y(n3678) );
  XOR2X1 U3480 ( .A(n3680), .B(N3000), .Y(n3677) );
  NOR4X1 U3481 ( .A(n3681), .B(n3682), .C(n3683), .D(n3684), .Y(n3668) );
  XNOR2X1 U3482 ( .A(N2985), .B(n3280), .Y(n3684) );
  MXI2X1 U3483 ( .A(N3733), .B(N2319), .S0(n3069), .Y(n3280) );
  XNOR2X1 U3484 ( .A(N2988), .B(n3685), .Y(n3683) );
  XNOR2X1 U3485 ( .A(N2984), .B(n3249), .Y(n3682) );
  MXI2X1 U3486 ( .A(N3732), .B(N2318), .S0(n3069), .Y(n3249) );
  NAND2X1 U3487 ( .A(n3686), .B(n3687), .Y(n3681) );
  XOR2X1 U3488 ( .A(n3688), .B(N2990), .Y(n3687) );
  XOR2X1 U3489 ( .A(n3689), .B(N2991), .Y(n3686) );
  NOR4X1 U3490 ( .A(n3690), .B(n3691), .C(n3692), .D(n3693), .Y(n3667) );
  XNOR2X1 U3491 ( .A(N2987), .B(n3694), .Y(n3693) );
  XNOR2X1 U3492 ( .A(N2997), .B(n3695), .Y(n3692) );
  XNOR2X1 U3493 ( .A(N2996), .B(n3696), .Y(n3691) );
  NAND2X1 U3494 ( .A(n3697), .B(n3698), .Y(n3690) );
  XOR2X1 U3495 ( .A(n3699), .B(N2999), .Y(n3698) );
  XOR2X1 U3496 ( .A(n3700), .B(N2986), .Y(n3697) );
  NOR4X1 U3497 ( .A(n3701), .B(n3702), .C(n3703), .D(n3704), .Y(n3666) );
  XNOR2X1 U3498 ( .A(N2992), .B(n3705), .Y(n3704) );
  XNOR2X1 U3499 ( .A(N2994), .B(n3706), .Y(n3703) );
  XNOR2X1 U3500 ( .A(N2993), .B(n3707), .Y(n3702) );
  NAND2X1 U3501 ( .A(n3708), .B(n3709), .Y(n3701) );
  XOR2X1 U3502 ( .A(n3710), .B(N2995), .Y(n3709) );
  XOR2X1 U3503 ( .A(n3711), .B(N2998), .Y(n3708) );
  OAI21XL U3504 ( .A0(n3332), .A1(n3483), .B0(n3524), .Y(n3664) );
  AOI2BB2X1 U3505 ( .B0(n3422), .B1(n3640), .A0N(n3342), .A1N(n3328), .Y(n3662) );
  CLKINVX1 U3506 ( .A(n3538), .Y(n3342) );
  NAND4X1 U3507 ( .A(n3713), .B(n3714), .C(n3715), .D(n3716), .Y(n3538) );
  NOR4X1 U3508 ( .A(n3717), .B(n3718), .C(n3719), .D(n3720), .Y(n3716) );
  XOR2X1 U3509 ( .A(N5164), .B(n3721), .Y(n3720) );
  XOR2X1 U3510 ( .A(N5166), .B(n3722), .Y(n3719) );
  XOR2X1 U3511 ( .A(N5165), .B(n3723), .Y(n3718) );
  NAND3X1 U3512 ( .A(n3724), .B(n3552), .C(n3725), .Y(n3717) );
  XNOR2X1 U3513 ( .A(n3726), .B(N5152), .Y(n3725) );
  CLKINVX1 U3514 ( .A(N5167), .Y(n3552) );
  XNOR2X1 U3515 ( .A(n3727), .B(N5163), .Y(n3724) );
  NOR4X1 U3516 ( .A(n3728), .B(n3729), .C(n3730), .D(n3731), .Y(n3715) );
  XNOR2X1 U3517 ( .A(N5148), .B(n3298), .Y(n3731) );
  MXI2X1 U3518 ( .A(N2319), .B(N3733), .S0(n3069), .Y(n3298) );
  XOR2X1 U3519 ( .A(N5151), .B(n3732), .Y(n3730) );
  XOR2X1 U3520 ( .A(N5147), .B(n3242), .Y(n3729) );
  CLKMX2X2 U3521 ( .A(N3732), .B(N2318), .S0(n3381), .Y(n3242) );
  NAND2X1 U3522 ( .A(n3733), .B(n3734), .Y(n3728) );
  XNOR2X1 U3523 ( .A(n3735), .B(N5153), .Y(n3734) );
  XNOR2X1 U3524 ( .A(n3736), .B(N5154), .Y(n3733) );
  NOR4X1 U3525 ( .A(n3737), .B(n3738), .C(n3739), .D(n3740), .Y(n3714) );
  XNOR2X1 U3526 ( .A(N5150), .B(n3741), .Y(n3740) );
  XOR2X1 U3527 ( .A(N5160), .B(n3742), .Y(n3739) );
  XOR2X1 U3528 ( .A(N5159), .B(n3743), .Y(n3738) );
  NAND2X1 U3529 ( .A(n3744), .B(n3745), .Y(n3737) );
  XNOR2X1 U3530 ( .A(n3746), .B(N5162), .Y(n3745) );
  XOR2X1 U3531 ( .A(n3747), .B(N5149), .Y(n3744) );
  NOR4X1 U3532 ( .A(n3748), .B(n3749), .C(n3750), .D(n3751), .Y(n3713) );
  XOR2X1 U3533 ( .A(N5155), .B(n3752), .Y(n3751) );
  XOR2X1 U3534 ( .A(N5157), .B(n3753), .Y(n3750) );
  XOR2X1 U3535 ( .A(N5156), .B(n3754), .Y(n3749) );
  NAND2X1 U3536 ( .A(n3755), .B(n3756), .Y(n3748) );
  XNOR2X1 U3537 ( .A(n3757), .B(N5158), .Y(n3756) );
  XNOR2X1 U3538 ( .A(n3758), .B(N5161), .Y(n3755) );
  MXI2X1 U3539 ( .A(n3759), .B(n3760), .S0(n3761), .Y(n3640) );
  NAND2BX1 U3540 ( .AN(n3762), .B(n3763), .Y(n3760) );
  AND2X1 U3541 ( .A(n3762), .B(n3763), .Y(n3522) );
  NOR3X1 U3542 ( .A(n3188), .B(n3426), .C(n3712), .Y(n3762) );
  NOR2X1 U3543 ( .A(n3645), .B(n3340), .Y(n3661) );
  CLKINVX1 U3544 ( .A(n3450), .Y(n3764) );
  MXI2X1 U3545 ( .A(n3765), .B(n3759), .S0(n3766), .Y(n3450) );
  MXI2X1 U3546 ( .A(n3338), .B(n2966), .S0(N3841), .Y(n3759) );
  AOI2BB1X1 U3547 ( .A0N(N3841), .A1N(n3348), .B0(n3763), .Y(n3765) );
  AND2X1 U3548 ( .A(N3841), .B(n3338), .Y(n3763) );
  CLKINVX1 U3549 ( .A(N6769), .Y(n3769) );
  OAI222XL U3550 ( .A0(n3771), .A1(n3767), .B0(n3772), .B1(n3768), .C0(n3770), 
        .C1(n3115), .Y(n1624) );
  CLKINVX1 U3551 ( .A(N6774), .Y(n3772) );
  OAI222XL U3552 ( .A0(n3773), .A1(n3767), .B0(n3774), .B1(n3768), .C0(n3770), 
        .C1(n2977), .Y(n1623) );
  CLKINVX1 U3553 ( .A(N6773), .Y(n3774) );
  OAI222XL U3554 ( .A0(n3775), .A1(n3767), .B0(n3776), .B1(n3768), .C0(n3770), 
        .C1(n2993), .Y(n1622) );
  CLKINVX1 U3555 ( .A(N6772), .Y(n3776) );
  CLKINVX1 U3556 ( .A(N6770), .Y(n3778) );
  OAI222XL U3557 ( .A0(n3779), .A1(n3767), .B0(n3768), .B1(n3780), .C0(n3770), 
        .C1(n2978), .Y(n1619) );
  CLKINVX1 U3558 ( .A(N6775), .Y(n3780) );
  NAND2X1 U3559 ( .A(n3181), .B(n3783), .Y(n3768) );
  NAND3X1 U3560 ( .A(n3782), .B(n3187), .C(n3781), .Y(n3767) );
  OAI21XL U3561 ( .A0(n3357), .A1(n3784), .B0(n3187), .Y(n3782) );
  MXI2X1 U3562 ( .A(n2984), .B(n3472), .S0(n3785), .Y(n1618) );
  CLKMX2X2 U3563 ( .A(pic_num[1]), .B(IM_Q[1]), .S0(n3785), .Y(n1617) );
  MXI2X1 U3564 ( .A(n2991), .B(n3474), .S0(n3785), .Y(n1616) );
  AND2X1 U3565 ( .A(n3786), .B(n3353), .Y(n3785) );
  MXI2X1 U3566 ( .A(n3789), .B(n3790), .S0(n4788), .Y(n1615) );
  OAI31XL U3567 ( .A0(n3791), .A1(pic_num[2]), .A2(n2991), .B0(n3790), .Y(
        n3789) );
  XOR2X1 U3568 ( .A(n2983), .B(n3792), .Y(n3791) );
  MXI2X1 U3569 ( .A(n3793), .B(n3794), .S0(n4787), .Y(n1614) );
  AOI21X1 U3570 ( .A0(n3795), .A1(n2981), .B0(n3796), .Y(n3794) );
  OR2X1 U3571 ( .A(n3792), .B(pic_num[2]), .Y(n3795) );
  NAND3X1 U3572 ( .A(n4788), .B(n3797), .C(n3790), .Y(n3793) );
  CLKINVX1 U3573 ( .A(n3796), .Y(n3790) );
  NAND4X1 U3574 ( .A(n3386), .B(n3186), .C(n3324), .D(n3798), .Y(n3796) );
  NOR4BBX1 U3575 ( .AN(n4705), .BN(n4706), .C(n3394), .D(n3799), .Y(n3324) );
  NAND4BX1 U3576 ( .AN(n3800), .B(n3801), .C(n3802), .D(n3803), .Y(n3394) );
  AND3X1 U3577 ( .A(n4697), .B(n4700), .C(n4699), .Y(n3803) );
  AND3X1 U3578 ( .A(n4691), .B(n4694), .C(n4692), .Y(n3802) );
  AND2X1 U3579 ( .A(n4690), .B(n4689), .Y(n3801) );
  NAND3BX1 U3580 ( .AN(n3804), .B(n4744), .C(n4745), .Y(n3800) );
  NOR2X1 U3581 ( .A(n3322), .B(n2980), .Y(n3186) );
  CLKINVX1 U3582 ( .A(n3392), .Y(n3322) );
  NOR2X1 U3583 ( .A(tick[2]), .B(tick[0]), .Y(n3392) );
  NOR2BX1 U3584 ( .AN(n3805), .B(n3354), .Y(n3386) );
  NAND3X1 U3585 ( .A(pic_num[1]), .B(n2984), .C(n3792), .Y(n3797) );
  NAND2X1 U3586 ( .A(pic_num[1]), .B(pic_num[0]), .Y(n3792) );
  MXI2X1 U3587 ( .A(n4800), .B(n3809), .S0(n3807), .Y(n1611) );
  MXI2X1 U3588 ( .A(n4801), .B(n3810), .S0(n3807), .Y(n1610) );
  MXI2X1 U3589 ( .A(n4802), .B(n3811), .S0(n3807), .Y(n1609) );
  MXI2X1 U3590 ( .A(n4803), .B(n3812), .S0(n3807), .Y(n1608) );
  MXI2X1 U3591 ( .A(n4804), .B(n3813), .S0(n3807), .Y(n1607) );
  MXI2X1 U3592 ( .A(n4805), .B(n3814), .S0(n3807), .Y(n1606) );
  MXI2X1 U3593 ( .A(n4806), .B(n3815), .S0(n3807), .Y(n1605) );
  MXI2X1 U3594 ( .A(n4807), .B(n3816), .S0(n3807), .Y(n1604) );
  MXI2X1 U3595 ( .A(n4790), .B(n3471), .S0(n3807), .Y(n1602) );
  MXI2X1 U3596 ( .A(n4791), .B(n3299), .S0(n3807), .Y(n1601) );
  MXI2X1 U3597 ( .A(n4792), .B(n3779), .S0(n3807), .Y(n1600) );
  MXI2X1 U3598 ( .A(n4793), .B(n3771), .S0(n3807), .Y(n1599) );
  MXI2X1 U3599 ( .A(n4794), .B(n3773), .S0(n3807), .Y(n1598) );
  MXI2X1 U3600 ( .A(n4795), .B(n3775), .S0(n3807), .Y(n1597) );
  AND2X1 U3601 ( .A(n3817), .B(n3818), .Y(n3364) );
  NOR2X1 U3602 ( .A(n3357), .B(n3784), .Y(n3786) );
  OAI2BB2XL U3603 ( .B0(n1420), .B1(n3819), .A0N(n3820), .A1N(n3821), .Y(n1593) );
  NAND4BX1 U3604 ( .AN(n3822), .B(n3823), .C(n3824), .D(n3825), .Y(n3821) );
  AOI222XL U3605 ( .A0(n3083), .A1(n3826), .B0(n3083), .B1(n3827), .C0(n3083), 
        .C1(n3828), .Y(n3825) );
  AOI22X1 U3606 ( .A0(n3083), .A1(n3829), .B0(n3083), .B1(n3830), .Y(n3824) );
  AOI22X1 U3607 ( .A0(n3083), .A1(n3831), .B0(n3083), .B1(n3832), .Y(n3823) );
  OAI211X1 U3608 ( .A0(n3833), .A1(n3002), .B0(n3834), .C0(n3835), .Y(n3822)
         );
  AO21X1 U3609 ( .A0(n3836), .A1(n3837), .B0(n3348), .Y(n3835) );
  AOI222XL U3610 ( .A0(n3083), .A1(n3838), .B0(n3083), .B1(n3839), .C0(n3083), 
        .C1(n3840), .Y(n3837) );
  AOI222XL U3611 ( .A0(n3083), .A1(n3841), .B0(n3083), .B1(n3842), .C0(n3083), 
        .C1(n3843), .Y(n3836) );
  AO21X1 U3612 ( .A0(n3844), .A1(n3845), .B0(n3467), .Y(n3834) );
  AOI222XL U3613 ( .A0(n3083), .A1(n3846), .B0(n3083), .B1(n3847), .C0(n3083), 
        .C1(n3848), .Y(n3845) );
  AOI222XL U3614 ( .A0(n3083), .A1(n3849), .B0(n3083), .B1(n3850), .C0(n3083), 
        .C1(n3851), .Y(n3844) );
  AOI222XL U3615 ( .A0(n3083), .A1(n3852), .B0(n3083), .B1(n3853), .C0(n3083), 
        .C1(n3854), .Y(n3833) );
  OAI2BB2XL U3616 ( .B0(n1419), .B1(n3819), .A0N(n3820), .A1N(n3855), .Y(n1592) );
  NAND4BX1 U3617 ( .AN(n3856), .B(n3857), .C(n3858), .D(n3859), .Y(n3855) );
  AOI222XL U3618 ( .A0(n3072), .A1(n3826), .B0(n3072), .B1(n3827), .C0(n3072), 
        .C1(n3828), .Y(n3859) );
  AOI22X1 U3619 ( .A0(n3072), .A1(n3829), .B0(n3072), .B1(n3830), .Y(n3858) );
  AOI22X1 U3620 ( .A0(n3072), .A1(n3831), .B0(n3072), .B1(n3832), .Y(n3857) );
  OAI211X1 U3621 ( .A0(n3860), .A1(n3002), .B0(n3861), .C0(n3862), .Y(n3856)
         );
  AO21X1 U3622 ( .A0(n3863), .A1(n3864), .B0(n3348), .Y(n3862) );
  AOI222XL U3623 ( .A0(n3072), .A1(n3838), .B0(n3072), .B1(n3839), .C0(n3072), 
        .C1(n3840), .Y(n3864) );
  AOI222XL U3624 ( .A0(n3072), .A1(n3841), .B0(n3072), .B1(n3842), .C0(n3072), 
        .C1(n3843), .Y(n3863) );
  AO21X1 U3625 ( .A0(n3865), .A1(n3866), .B0(n3467), .Y(n3861) );
  AOI222XL U3626 ( .A0(n3072), .A1(n3846), .B0(n3072), .B1(n3847), .C0(n3072), 
        .C1(n3848), .Y(n3866) );
  AOI222XL U3627 ( .A0(n3072), .A1(n3849), .B0(n3072), .B1(n3850), .C0(n3072), 
        .C1(n3851), .Y(n3865) );
  AOI222XL U3628 ( .A0(n3072), .A1(n3852), .B0(n3072), .B1(n3853), .C0(n3072), 
        .C1(n3854), .Y(n3860) );
  OAI2BB2XL U3629 ( .B0(n1418), .B1(n3819), .A0N(n3820), .A1N(n3867), .Y(n1591) );
  NAND4BX1 U3630 ( .AN(n3868), .B(n3869), .C(n3870), .D(n3871), .Y(n3867) );
  AOI222XL U3631 ( .A0(n3071), .A1(n3826), .B0(n3071), .B1(n3827), .C0(n3071), 
        .C1(n3828), .Y(n3871) );
  AOI22X1 U3632 ( .A0(n3071), .A1(n3829), .B0(n3071), .B1(n3830), .Y(n3870) );
  AOI22X1 U3633 ( .A0(n3071), .A1(n3831), .B0(n3071), .B1(n3832), .Y(n3869) );
  OAI211X1 U3634 ( .A0(n3872), .A1(n3002), .B0(n3873), .C0(n3874), .Y(n3868)
         );
  AO21X1 U3635 ( .A0(n3875), .A1(n3876), .B0(n3348), .Y(n3874) );
  AOI222XL U3636 ( .A0(n3071), .A1(n3838), .B0(n3071), .B1(n3839), .C0(n3071), 
        .C1(n3840), .Y(n3876) );
  AOI222XL U3637 ( .A0(n3071), .A1(n3841), .B0(n3071), .B1(n3842), .C0(n3071), 
        .C1(n3843), .Y(n3875) );
  AO21X1 U3638 ( .A0(n3877), .A1(n3878), .B0(n3467), .Y(n3873) );
  AOI222XL U3639 ( .A0(n3071), .A1(n3846), .B0(n3071), .B1(n3847), .C0(n3071), 
        .C1(n3848), .Y(n3878) );
  AOI222XL U3640 ( .A0(n3071), .A1(n3849), .B0(n3071), .B1(n3850), .C0(n3071), 
        .C1(n3851), .Y(n3877) );
  AOI222XL U3641 ( .A0(n3071), .A1(n3852), .B0(n3071), .B1(n3853), .C0(n3071), 
        .C1(n3854), .Y(n3872) );
  OAI2BB2XL U3642 ( .B0(n1417), .B1(n3819), .A0N(n3820), .A1N(n3879), .Y(n1590) );
  NAND4BX1 U3643 ( .AN(n3880), .B(n3881), .C(n3882), .D(n3883), .Y(n3879) );
  AOI222XL U3644 ( .A0(n3016), .A1(n3826), .B0(n2982), .B1(n3827), .C0(n2982), 
        .C1(n3828), .Y(n3883) );
  AOI22X1 U3645 ( .A0(n3016), .A1(n3831), .B0(n2982), .B1(n3832), .Y(n3881) );
  OAI211X1 U3646 ( .A0(n3884), .A1(n3002), .B0(n3885), .C0(n3886), .Y(n3880)
         );
  AO21X1 U3647 ( .A0(n3887), .A1(n3888), .B0(n3348), .Y(n3886) );
  AOI222XL U3648 ( .A0(N6436), .A1(n3838), .B0(N6410), .B1(n3839), .C0(N6383), 
        .C1(n3840), .Y(n3888) );
  AOI222XL U3649 ( .A0(N6302), .A1(n3841), .B0(N6329), .B1(n3842), .C0(N6356), 
        .C1(n3843), .Y(n3887) );
  AO21X1 U3650 ( .A0(n3889), .A1(n3890), .B0(n3467), .Y(n3885) );
  AOI222XL U3651 ( .A0(N6195), .A1(n3846), .B0(N6169), .B1(n3847), .C0(N6142), 
        .C1(n3848), .Y(n3890) );
  AOI222XL U3652 ( .A0(N6061), .A1(n3849), .B0(N6088), .B1(n3850), .C0(N6115), 
        .C1(n3851), .Y(n3889) );
  AOI222XL U3653 ( .A0(N5892), .A1(n3852), .B0(N5919), .B1(n3853), .C0(N5945), 
        .C1(n3854), .Y(n3884) );
  OAI2BB2XL U3654 ( .B0(n1416), .B1(n3819), .A0N(n3820), .A1N(n3891), .Y(n1589) );
  NAND4BX1 U3655 ( .AN(n3892), .B(n3893), .C(n3894), .D(n3895), .Y(n3891) );
  AOI222XL U3656 ( .A0(n3075), .A1(n3826), .B0(N6024), .B1(n3827), .C0(N5852), 
        .C1(n3828), .Y(n3895) );
  AOI22X1 U3657 ( .A0(n3075), .A1(n3831), .B0(N6005), .B1(n3832), .Y(n3893) );
  OAI211X1 U3658 ( .A0(n3896), .A1(n3002), .B0(n3897), .C0(n3898), .Y(n3892)
         );
  AO21X1 U3659 ( .A0(n3899), .A1(n3900), .B0(n3348), .Y(n3898) );
  AOI222XL U3660 ( .A0(N6437), .A1(n3838), .B0(N6411), .B1(n3839), .C0(N6384), 
        .C1(n3840), .Y(n3900) );
  AOI222XL U3661 ( .A0(N6303), .A1(n3841), .B0(N6330), .B1(n3842), .C0(N6357), 
        .C1(n3843), .Y(n3899) );
  AO21X1 U3662 ( .A0(n3901), .A1(n3902), .B0(n3467), .Y(n3897) );
  AOI222XL U3663 ( .A0(N6196), .A1(n3846), .B0(N6170), .B1(n3847), .C0(N6143), 
        .C1(n3848), .Y(n3902) );
  AOI222XL U3664 ( .A0(N6062), .A1(n3849), .B0(N6089), .B1(n3850), .C0(N6116), 
        .C1(n3851), .Y(n3901) );
  AOI222XL U3665 ( .A0(N5893), .A1(n3852), .B0(N5920), .B1(n3853), .C0(N5946), 
        .C1(n3854), .Y(n3896) );
  OAI2BB2XL U3666 ( .B0(n1415), .B1(n3819), .A0N(n3820), .A1N(n3903), .Y(n1588) );
  NAND4BX1 U3667 ( .AN(n3904), .B(n3905), .C(n3906), .D(n3907), .Y(n3903) );
  AOI222XL U3668 ( .A0(n3081), .A1(n3826), .B0(N6025), .B1(n3827), .C0(N5853), 
        .C1(n3828), .Y(n3907) );
  AOI22X1 U3669 ( .A0(n3080), .A1(n3831), .B0(N6006), .B1(n3832), .Y(n3905) );
  OAI211X1 U3670 ( .A0(n3908), .A1(n3002), .B0(n3909), .C0(n3910), .Y(n3904)
         );
  AO21X1 U3671 ( .A0(n3911), .A1(n3912), .B0(n3348), .Y(n3910) );
  AOI222XL U3672 ( .A0(N6438), .A1(n3838), .B0(N6412), .B1(n3839), .C0(N6385), 
        .C1(n3840), .Y(n3912) );
  AOI222XL U3673 ( .A0(N6304), .A1(n3841), .B0(N6331), .B1(n3842), .C0(N6358), 
        .C1(n3843), .Y(n3911) );
  AO21X1 U3674 ( .A0(n3913), .A1(n3914), .B0(n3467), .Y(n3909) );
  AOI222XL U3675 ( .A0(N6197), .A1(n3846), .B0(N6171), .B1(n3847), .C0(N6144), 
        .C1(n3848), .Y(n3914) );
  AOI222XL U3676 ( .A0(N6063), .A1(n3849), .B0(N6090), .B1(n3850), .C0(N6117), 
        .C1(n3851), .Y(n3913) );
  AOI222XL U3677 ( .A0(N5894), .A1(n3852), .B0(N5921), .B1(n3853), .C0(N5947), 
        .C1(n3854), .Y(n3908) );
  OAI2BB2XL U3678 ( .B0(n1414), .B1(n3819), .A0N(n3820), .A1N(n3915), .Y(n1587) );
  NAND4BX1 U3679 ( .AN(n3916), .B(n3917), .C(n3918), .D(n3919), .Y(n3915) );
  AOI222XL U3680 ( .A0(n3077), .A1(n3826), .B0(N6026), .B1(n3827), .C0(N5854), 
        .C1(n3828), .Y(n3919) );
  AOI22X1 U3681 ( .A0(N6017), .A1(n3831), .B0(N6007), .B1(n3832), .Y(n3917) );
  OAI211X1 U3682 ( .A0(n3920), .A1(n3002), .B0(n3921), .C0(n3922), .Y(n3916)
         );
  AO21X1 U3683 ( .A0(n3923), .A1(n3924), .B0(n3348), .Y(n3922) );
  AOI222XL U3684 ( .A0(N6439), .A1(n3838), .B0(N6413), .B1(n3839), .C0(N6386), 
        .C1(n3840), .Y(n3924) );
  AOI222XL U3685 ( .A0(N6305), .A1(n3841), .B0(N6332), .B1(n3842), .C0(N6359), 
        .C1(n3843), .Y(n3923) );
  AO21X1 U3686 ( .A0(n3925), .A1(n3926), .B0(n3467), .Y(n3921) );
  AOI222XL U3687 ( .A0(N6198), .A1(n3846), .B0(N6172), .B1(n3847), .C0(N6145), 
        .C1(n3848), .Y(n3926) );
  AOI222XL U3688 ( .A0(N6064), .A1(n3849), .B0(N6091), .B1(n3850), .C0(N6118), 
        .C1(n3851), .Y(n3925) );
  AOI222XL U3689 ( .A0(N5895), .A1(n3852), .B0(N5922), .B1(n3853), .C0(N5948), 
        .C1(n3854), .Y(n3920) );
  OAI2BB2XL U3690 ( .B0(n1413), .B1(n3819), .A0N(n3820), .A1N(n3927), .Y(n1586) );
  NAND4BX1 U3691 ( .AN(n3928), .B(n3929), .C(n3930), .D(n3931), .Y(n3927) );
  AOI222XL U3692 ( .A0(n3079), .A1(n3826), .B0(N6027), .B1(n3827), .C0(N5855), 
        .C1(n3828), .Y(n3931) );
  AOI22X1 U3693 ( .A0(N6018), .A1(n3831), .B0(N6008), .B1(n3832), .Y(n3929) );
  OAI211X1 U3694 ( .A0(n3932), .A1(n3002), .B0(n3933), .C0(n3934), .Y(n3928)
         );
  AO21X1 U3695 ( .A0(n3935), .A1(n3936), .B0(n3348), .Y(n3934) );
  AOI222XL U3696 ( .A0(N6440), .A1(n3838), .B0(N6414), .B1(n3839), .C0(N6387), 
        .C1(n3840), .Y(n3936) );
  AOI222XL U3697 ( .A0(N6306), .A1(n3841), .B0(N6333), .B1(n3842), .C0(N6360), 
        .C1(n3843), .Y(n3935) );
  AO21X1 U3698 ( .A0(n3937), .A1(n3938), .B0(n3467), .Y(n3933) );
  AOI222XL U3699 ( .A0(N6199), .A1(n3846), .B0(N6173), .B1(n3847), .C0(N6146), 
        .C1(n3848), .Y(n3938) );
  AOI222XL U3700 ( .A0(N6065), .A1(n3849), .B0(N6092), .B1(n3850), .C0(N6119), 
        .C1(n3851), .Y(n3937) );
  AOI222XL U3701 ( .A0(N5896), .A1(n3852), .B0(N5923), .B1(n3853), .C0(N5949), 
        .C1(n3854), .Y(n3932) );
  OAI2BB2XL U3702 ( .B0(n1412), .B1(n3819), .A0N(n3820), .A1N(n3939), .Y(n1585) );
  NAND4BX1 U3703 ( .AN(n3940), .B(n3941), .C(n3942), .D(n3943), .Y(n3939) );
  AOI222XL U3704 ( .A0(n3073), .A1(n3826), .B0(N6028), .B1(n3827), .C0(N5856), 
        .C1(n3828), .Y(n3943) );
  AOI222XL U3705 ( .A0(n3338), .A1(n3850), .B0(n3842), .B1(n3945), .C0(n3946), 
        .C1(n3853), .Y(n3944) );
  AOI222XL U3706 ( .A0(n3338), .A1(n3851), .B0(n3843), .B1(n3945), .C0(n3854), 
        .C1(n3946), .Y(n3953) );
  AOI22X1 U3707 ( .A0(N6019), .A1(n3831), .B0(N6009), .B1(n3832), .Y(n3941) );
  OAI211X1 U3708 ( .A0(n3956), .A1(n3002), .B0(n3957), .C0(n3958), .Y(n3940)
         );
  AO21X1 U3709 ( .A0(n3959), .A1(n3960), .B0(n3348), .Y(n3958) );
  AOI222XL U3710 ( .A0(N6441), .A1(n3838), .B0(N6415), .B1(n3839), .C0(N6388), 
        .C1(n3840), .Y(n3960) );
  NAND2X1 U3711 ( .A(n3961), .B(n3962), .Y(n3954) );
  CLKINVX1 U3712 ( .A(n3965), .Y(n3964) );
  NAND2X1 U3713 ( .A(n3966), .B(n2978), .Y(n3963) );
  OAI31XL U3714 ( .A0(N6391), .A1(sec[3]), .A2(N6392), .B0(sec[4]), .Y(n3966)
         );
  AOI222XL U3715 ( .A0(N6307), .A1(n3841), .B0(N6334), .B1(n3842), .C0(N6361), 
        .C1(n3843), .Y(n3959) );
  NAND2X1 U3716 ( .A(n3965), .B(n3968), .Y(n3962) );
  NAND4X1 U3717 ( .A(N6391), .B(N6392), .C(sec[3]), .D(sec[4]), .Y(n3968) );
  NAND2X1 U3718 ( .A(n3965), .B(n3969), .Y(n3967) );
  OAI21XL U3719 ( .A0(sec[3]), .A1(N6392), .B0(sec[4]), .Y(n3969) );
  NAND3X1 U3720 ( .A(n3970), .B(n2977), .C(n3965), .Y(n3948) );
  NOR2X1 U3721 ( .A(sec[5]), .B(sec[6]), .Y(n3965) );
  OAI21XL U3722 ( .A0(N6392), .A1(N6391), .B0(sec[3]), .Y(n3970) );
  AO21X1 U3723 ( .A0(n3971), .A1(n3972), .B0(n3467), .Y(n3957) );
  AOI222XL U3724 ( .A0(N6200), .A1(n3846), .B0(N6174), .B1(n3847), .C0(N6147), 
        .C1(n3848), .Y(n3972) );
  NAND2X1 U3725 ( .A(n3973), .B(n3974), .Y(n3955) );
  CLKINVX1 U3726 ( .A(n3976), .Y(n3973) );
  AOI31X1 U3727 ( .A0(n4866), .A1(n4868), .A2(n4865), .B0(n3977), .Y(n3976) );
  NAND2X1 U3728 ( .A(n4865), .B(n3978), .Y(n3975) );
  OAI31XL U3729 ( .A0(n3979), .A1(N6150), .A2(n3980), .B0(min[4]), .Y(n3978)
         );
  AOI222XL U3730 ( .A0(N6066), .A1(n3849), .B0(N6093), .B1(n3850), .C0(N6120), 
        .C1(n3851), .Y(n3971) );
  OAI21XL U3731 ( .A0(n4869), .A1(n3982), .B0(n3977), .Y(n3974) );
  NAND2X1 U3732 ( .A(n3977), .B(n3983), .Y(n3981) );
  OAI21XL U3733 ( .A0(n3980), .A1(n3979), .B0(min[4]), .Y(n3983) );
  NAND3X1 U3734 ( .A(n4866), .B(n3984), .C(n3977), .Y(n3947) );
  AND2X1 U3735 ( .A(n4864), .B(n4865), .Y(n3977) );
  OAI21XL U3736 ( .A0(N6150), .A1(n3979), .B0(n3980), .Y(n3984) );
  AOI222XL U3737 ( .A0(N5897), .A1(n3852), .B0(N5924), .B1(n3853), .C0(N5950), 
        .C1(n3854), .Y(n3956) );
  AO21X1 U3738 ( .A0(n4863), .A1(n4862), .B0(n4861), .Y(n3985) );
  NAND4X1 U3739 ( .A(n4859), .B(n4860), .C(n4861), .D(n3986), .Y(n3951) );
  AO21X1 U3740 ( .A0(n4863), .A1(n4858), .B0(n4862), .Y(n3986) );
  NAND2X1 U3741 ( .A(n3475), .B(n3365), .Y(n3784) );
  NOR2X1 U3742 ( .A(n2964), .B(n3989), .Y(n3952) );
  OAI22XL U3743 ( .A0(n2110), .A1(n3991), .B0(n3470), .B1(n3992), .Y(n1584) );
  OAI22XL U3744 ( .A0(n2111), .A1(n3991), .B0(n3471), .B1(n3992), .Y(n1583) );
  OAI22XL U3745 ( .A0(n2112), .A1(n3991), .B0(n3299), .B1(n3992), .Y(n1582) );
  OAI22XL U3746 ( .A0(n2113), .A1(n3991), .B0(n3779), .B1(n3992), .Y(n1581) );
  OAI22XL U3747 ( .A0(n2114), .A1(n3991), .B0(n3771), .B1(n3992), .Y(n1580) );
  OAI22XL U3748 ( .A0(n2115), .A1(n3991), .B0(n3773), .B1(n3992), .Y(n1579) );
  OAI22XL U3749 ( .A0(n2116), .A1(n3991), .B0(n3775), .B1(n3992), .Y(n1578) );
  OAI22XL U3750 ( .A0(n2117), .A1(n3991), .B0(n3472), .B1(n3992), .Y(n1577) );
  OAI22XL U3751 ( .A0(n2118), .A1(n3991), .B0(n3992), .B1(n3993), .Y(n1576) );
  OAI22XL U3752 ( .A0(n2119), .A1(n3991), .B0(n3992), .B1(n3994), .Y(n1575) );
  OAI22XL U3753 ( .A0(n2120), .A1(n3991), .B0(n3992), .B1(n3995), .Y(n1574) );
  OAI22XL U3754 ( .A0(n2121), .A1(n3991), .B0(n3992), .B1(n3996), .Y(n1573) );
  OAI22XL U3755 ( .A0(n2122), .A1(n3991), .B0(n3473), .B1(n3992), .Y(n1572) );
  OAI22XL U3756 ( .A0(n2123), .A1(n3991), .B0(n3806), .B1(n3992), .Y(n1571) );
  OAI22XL U3757 ( .A0(n2124), .A1(n3991), .B0(n3808), .B1(n3992), .Y(n1570) );
  OAI22XL U3758 ( .A0(n2125), .A1(n3991), .B0(n3809), .B1(n3992), .Y(n1569) );
  OAI22XL U3759 ( .A0(n2126), .A1(n3991), .B0(n3810), .B1(n3992), .Y(n1568) );
  OAI22XL U3760 ( .A0(n2127), .A1(n3991), .B0(n3811), .B1(n3992), .Y(n1567) );
  OAI22XL U3761 ( .A0(n2128), .A1(n3991), .B0(n3812), .B1(n3992), .Y(n1566) );
  OAI22XL U3762 ( .A0(n2129), .A1(n3991), .B0(n3813), .B1(n3992), .Y(n1565) );
  OAI22XL U3763 ( .A0(n2130), .A1(n3991), .B0(n3814), .B1(n3992), .Y(n1564) );
  OAI22XL U3764 ( .A0(n2131), .A1(n3991), .B0(n3815), .B1(n3992), .Y(n1563) );
  OAI22XL U3765 ( .A0(n2132), .A1(n3991), .B0(n3816), .B1(n3992), .Y(n1562) );
  OAI22XL U3766 ( .A0(n2133), .A1(n3991), .B0(n3474), .B1(n3992), .Y(n1561) );
  MXI2X1 U3767 ( .A(n3998), .B(n3999), .S0(n3946), .Y(n3997) );
  NAND3X1 U3768 ( .A(n3367), .B(n4000), .C(n3531), .Y(n3999) );
  OAI21XL U3769 ( .A0(N444), .A1(n3451), .B0(n3379), .Y(n4000) );
  NAND2X1 U3770 ( .A(n3989), .B(n4001), .Y(n3998) );
  OR2X1 U3771 ( .A(n3989), .B(n3458), .Y(n4003) );
  NOR2X1 U3772 ( .A(n4004), .B(n4854), .Y(n3989) );
  OAI31XL U3773 ( .A0(n4005), .A1(n3343), .A2(n3950), .B0(n3367), .Y(n4002) );
  OAI21XL U3774 ( .A0(n3451), .A1(n3478), .B0(n3201), .Y(n4005) );
  MXI2X1 U3775 ( .A(n4819), .B(n3993), .S0(n3070), .Y(n1512) );
  CLKINVX1 U3776 ( .A(IM_Q[23]), .Y(n3993) );
  MXI2X1 U3777 ( .A(n4820), .B(n3994), .S0(n3070), .Y(n1511) );
  MXI2X1 U3778 ( .A(n4821), .B(n3995), .S0(n3070), .Y(n1510) );
  MXI2X1 U3779 ( .A(n4822), .B(n3996), .S0(n3070), .Y(n1509) );
  MXI2X1 U3780 ( .A(n4824), .B(n3806), .S0(n3070), .Y(n1508) );
  MXI2X1 U3781 ( .A(n4825), .B(n3808), .S0(n3070), .Y(n1507) );
  MXI2X1 U3782 ( .A(n4826), .B(n3809), .S0(n3070), .Y(n1506) );
  MXI2X1 U3783 ( .A(n4827), .B(n3810), .S0(n3070), .Y(n1505) );
  MXI2X1 U3784 ( .A(n4828), .B(n3811), .S0(n3070), .Y(n1504) );
  MXI2X1 U3785 ( .A(n4829), .B(n3812), .S0(n3070), .Y(n1503) );
  MXI2X1 U3786 ( .A(n4830), .B(n3813), .S0(n3070), .Y(n1502) );
  MXI2X1 U3787 ( .A(n4831), .B(n3814), .S0(n3070), .Y(n1501) );
  MXI2X1 U3788 ( .A(n4832), .B(n3815), .S0(n3070), .Y(n1500) );
  MXI2X1 U3789 ( .A(n4833), .B(n3816), .S0(n3070), .Y(n1499) );
  MXI2X1 U3790 ( .A(n4811), .B(n3470), .S0(n3070), .Y(n1498) );
  MXI2X1 U3791 ( .A(n4778), .B(n3471), .S0(n3070), .Y(n1497) );
  MXI2X1 U3792 ( .A(n4779), .B(n3299), .S0(n3070), .Y(n1496) );
  MXI2X1 U3793 ( .A(n4780), .B(n3779), .S0(n3070), .Y(n1495) );
  MXI2X1 U3794 ( .A(n4781), .B(n3771), .S0(n3070), .Y(n1494) );
  MXI2X1 U3795 ( .A(n4782), .B(n3773), .S0(n3070), .Y(n1493) );
  MXI2X1 U3796 ( .A(n4783), .B(n3775), .S0(n3070), .Y(n1492) );
  MXI2X1 U3797 ( .A(n4784), .B(n3472), .S0(n3070), .Y(n1491) );
  MXI2X1 U3798 ( .A(n4785), .B(n3473), .S0(n3070), .Y(n1490) );
  MXI2X1 U3799 ( .A(n4786), .B(n3474), .S0(n3070), .Y(n1489) );
  NOR2BX1 U3800 ( .AN(n4007), .B(n2996), .Y(n4009) );
  NAND4BX1 U3801 ( .AN(n4010), .B(n4011), .C(n4012), .D(n4013), .Y(n1488) );
  AOI221XL U3802 ( .A0(N3165), .A1(n4014), .B0(n3410), .B1(n4015), .C0(n4016), 
        .Y(n4013) );
  OAI2BB2XL U3803 ( .B0(n4017), .B1(n3347), .A0N(n4018), .A1N(N250), .Y(n4015)
         );
  NOR4X1 U3804 ( .A(n4019), .B(n4020), .C(n4021), .D(n4022), .Y(n4017) );
  OAI22XL U3805 ( .A0(n4823), .A1(n4023), .B0(n4785), .B1(n3950), .Y(n4022) );
  OAI22XL U3806 ( .A0(n4766), .A1(n4024), .B0(n3949), .B1(n4025), .Y(n4021) );
  OAI22XL U3807 ( .A0(n4752), .A1(n3467), .B0(n2996), .B1(n4026), .Y(n4020) );
  OAI2BB2XL U3808 ( .B0(n2122), .B1(n4027), .A0N(N4272), .A1N(n4028), .Y(n4019) );
  OA22X1 U3809 ( .A0(n4029), .A1(n4823), .B0(n4030), .B1(n3440), .Y(n4012) );
  AOI222XL U3810 ( .A0(N2183), .A1(n4031), .B0(IM_Q[1]), .B1(n4032), .C0(N250), 
        .C1(n4018), .Y(n4030) );
  OA22X1 U3811 ( .A0(n4025), .A1(n4033), .B0(n4026), .B1(n4034), .Y(n4011) );
  CLKINVX1 U3812 ( .A(N3689), .Y(n4026) );
  CLKINVX1 U3813 ( .A(N3664), .Y(n4025) );
  OAI22XL U3814 ( .A0(n4752), .A1(n4035), .B0(n4785), .B1(n4036), .Y(n4010) );
  NAND4BX1 U3815 ( .AN(n4037), .B(n4038), .C(n4039), .D(n4040), .Y(n1487) );
  AOI221XL U3816 ( .A0(N3166), .A1(n4014), .B0(n3410), .B1(n4041), .C0(n4016), 
        .Y(n4040) );
  OAI2BB2XL U3817 ( .B0(n4042), .B1(n3347), .A0N(n4018), .A1N(N249), .Y(n4041)
         );
  NOR4X1 U3818 ( .A(n4043), .B(n4044), .C(n4045), .D(n4046), .Y(n4042) );
  OAI22XL U3819 ( .A0(n4818), .A1(n4023), .B0(n4784), .B1(n3950), .Y(n4046) );
  OAI22XL U3820 ( .A0(n4761), .A1(n4024), .B0(n3949), .B1(n4047), .Y(n4045) );
  OAI22XL U3821 ( .A0(n4751), .A1(n3467), .B0(n2996), .B1(n4048), .Y(n4044) );
  OAI2BB2XL U3822 ( .B0(n2117), .B1(n4027), .A0N(N4273), .A1N(n4028), .Y(n4043) );
  OA22X1 U3823 ( .A0(n4029), .A1(n4818), .B0(n4049), .B1(n3440), .Y(n4039) );
  AOI222XL U3824 ( .A0(N2184), .A1(n4031), .B0(IM_Q[2]), .B1(n4032), .C0(N249), 
        .C1(n4018), .Y(n4049) );
  OA22X1 U3825 ( .A0(n4033), .A1(n4047), .B0(n4034), .B1(n4048), .Y(n4038) );
  CLKINVX1 U3826 ( .A(N3690), .Y(n4048) );
  CLKINVX1 U3827 ( .A(N3665), .Y(n4047) );
  OAI22XL U3828 ( .A0(n4751), .A1(n4035), .B0(n4784), .B1(n4036), .Y(n4037) );
  NAND4BX1 U3829 ( .AN(n4050), .B(n4051), .C(n4052), .D(n4053), .Y(n1486) );
  AOI221XL U3830 ( .A0(N3167), .A1(n4014), .B0(n3410), .B1(n4054), .C0(n4016), 
        .Y(n4053) );
  OAI2BB2XL U3831 ( .B0(n4055), .B1(n3347), .A0N(n4018), .A1N(N248), .Y(n4054)
         );
  NOR4X1 U3832 ( .A(n4056), .B(n4057), .C(n4058), .D(n4059), .Y(n4055) );
  OAI22XL U3833 ( .A0(n4817), .A1(n4023), .B0(n4783), .B1(n3950), .Y(n4059) );
  OAI22XL U3834 ( .A0(n4760), .A1(n4024), .B0(n3949), .B1(n4060), .Y(n4058) );
  OAI22XL U3835 ( .A0(n4750), .A1(n3467), .B0(n2996), .B1(n4061), .Y(n4057) );
  OAI2BB2XL U3836 ( .B0(n2116), .B1(n4027), .A0N(N4274), .A1N(n4028), .Y(n4056) );
  OA22X1 U3837 ( .A0(n4029), .A1(n4817), .B0(n4062), .B1(n3440), .Y(n4052) );
  AOI222XL U3838 ( .A0(N2185), .A1(n4031), .B0(IM_Q[3]), .B1(n4032), .C0(N248), 
        .C1(n4018), .Y(n4062) );
  OA22X1 U3839 ( .A0(n4033), .A1(n4060), .B0(n4034), .B1(n4061), .Y(n4051) );
  CLKINVX1 U3840 ( .A(N3691), .Y(n4061) );
  CLKINVX1 U3841 ( .A(N3666), .Y(n4060) );
  OAI22XL U3842 ( .A0(n4750), .A1(n4035), .B0(n4783), .B1(n4036), .Y(n4050) );
  NAND4BX1 U3843 ( .AN(n4063), .B(n4064), .C(n4065), .D(n4066), .Y(n1485) );
  AOI221XL U3844 ( .A0(N3168), .A1(n4014), .B0(n3410), .B1(n4067), .C0(n4016), 
        .Y(n4066) );
  OAI2BB2XL U3845 ( .B0(n4068), .B1(n3347), .A0N(n4018), .A1N(N247), .Y(n4067)
         );
  NOR4X1 U3846 ( .A(n4069), .B(n4070), .C(n4071), .D(n4072), .Y(n4068) );
  OAI22XL U3847 ( .A0(n4816), .A1(n4023), .B0(n4782), .B1(n3950), .Y(n4072) );
  OAI22XL U3848 ( .A0(n4759), .A1(n4024), .B0(n3949), .B1(n4073), .Y(n4071) );
  OAI22XL U3849 ( .A0(n4749), .A1(n3467), .B0(n2996), .B1(n4074), .Y(n4070) );
  OAI2BB2XL U3850 ( .B0(n2115), .B1(n4027), .A0N(N4275), .A1N(n4028), .Y(n4069) );
  OA22X1 U3851 ( .A0(n4029), .A1(n4816), .B0(n4075), .B1(n3440), .Y(n4065) );
  AOI222XL U3852 ( .A0(N2186), .A1(n4031), .B0(IM_Q[4]), .B1(n4032), .C0(N247), 
        .C1(n4018), .Y(n4075) );
  OA22X1 U3853 ( .A0(n4033), .A1(n4073), .B0(n4034), .B1(n4074), .Y(n4064) );
  CLKINVX1 U3854 ( .A(N3692), .Y(n4074) );
  CLKINVX1 U3855 ( .A(N3667), .Y(n4073) );
  OAI22XL U3856 ( .A0(n4749), .A1(n4035), .B0(n4782), .B1(n4036), .Y(n4063) );
  NAND4BX1 U3857 ( .AN(n4076), .B(n4077), .C(n4078), .D(n4079), .Y(n1484) );
  AOI221XL U3858 ( .A0(N3169), .A1(n4014), .B0(n3410), .B1(n4080), .C0(n4016), 
        .Y(n4079) );
  OAI2BB2XL U3859 ( .B0(n4081), .B1(n3347), .A0N(n4018), .A1N(N246), .Y(n4080)
         );
  NOR4X1 U3860 ( .A(n4082), .B(n4083), .C(n4084), .D(n4085), .Y(n4081) );
  OAI22XL U3861 ( .A0(n4815), .A1(n4023), .B0(n4781), .B1(n3950), .Y(n4085) );
  OAI22XL U3862 ( .A0(n4758), .A1(n4024), .B0(n3949), .B1(n4086), .Y(n4084) );
  OAI22XL U3863 ( .A0(n4748), .A1(n3467), .B0(n2996), .B1(n4087), .Y(n4083) );
  OAI2BB2XL U3864 ( .B0(n2114), .B1(n4027), .A0N(N4276), .A1N(n4028), .Y(n4082) );
  OA22X1 U3865 ( .A0(n4029), .A1(n4815), .B0(n4088), .B1(n3440), .Y(n4078) );
  AOI222XL U3866 ( .A0(N2187), .A1(n4031), .B0(IM_Q[5]), .B1(n4032), .C0(N246), 
        .C1(n4018), .Y(n4088) );
  OA22X1 U3867 ( .A0(n4033), .A1(n4086), .B0(n4034), .B1(n4087), .Y(n4077) );
  CLKINVX1 U3868 ( .A(N3693), .Y(n4087) );
  CLKINVX1 U3869 ( .A(N3668), .Y(n4086) );
  OAI22XL U3870 ( .A0(n4748), .A1(n4035), .B0(n4781), .B1(n4036), .Y(n4076) );
  NAND4BX1 U3871 ( .AN(n4089), .B(n4090), .C(n4091), .D(n4092), .Y(n1483) );
  AOI221XL U3872 ( .A0(N3170), .A1(n4014), .B0(n3410), .B1(n4093), .C0(n4016), 
        .Y(n4092) );
  OAI2BB2XL U3873 ( .B0(n4094), .B1(n3347), .A0N(n4018), .A1N(N245), .Y(n4093)
         );
  NOR4X1 U3874 ( .A(n4095), .B(n4096), .C(n4097), .D(n4098), .Y(n4094) );
  OAI22XL U3875 ( .A0(n4814), .A1(n4023), .B0(n4780), .B1(n3950), .Y(n4098) );
  OAI22XL U3876 ( .A0(n4757), .A1(n4024), .B0(n3949), .B1(n4099), .Y(n4097) );
  OAI22XL U3877 ( .A0(n4747), .A1(n3467), .B0(n2996), .B1(n4100), .Y(n4096) );
  OAI2BB2XL U3878 ( .B0(n2113), .B1(n4027), .A0N(N4277), .A1N(n4028), .Y(n4095) );
  OA22X1 U3879 ( .A0(n4029), .A1(n4814), .B0(n4101), .B1(n3440), .Y(n4091) );
  AOI222XL U3880 ( .A0(N2188), .A1(n4031), .B0(IM_Q[6]), .B1(n4032), .C0(N245), 
        .C1(n4018), .Y(n4101) );
  OA22X1 U3881 ( .A0(n4033), .A1(n4099), .B0(n4034), .B1(n4100), .Y(n4090) );
  CLKINVX1 U3882 ( .A(N3694), .Y(n4100) );
  CLKINVX1 U3883 ( .A(N3669), .Y(n4099) );
  OAI22XL U3884 ( .A0(n4747), .A1(n4035), .B0(n4780), .B1(n4036), .Y(n4089) );
  NAND4BX1 U3885 ( .AN(n4102), .B(n4103), .C(n4104), .D(n4105), .Y(n1482) );
  AOI221XL U3886 ( .A0(N3171), .A1(n4014), .B0(n3410), .B1(n4106), .C0(n4016), 
        .Y(n4105) );
  OAI2BB2XL U3887 ( .B0(n4107), .B1(n3347), .A0N(n4018), .A1N(N244), .Y(n4106)
         );
  NOR4X1 U3888 ( .A(n4108), .B(n4109), .C(n4110), .D(n4111), .Y(n4107) );
  OAI22XL U3889 ( .A0(n4813), .A1(n4023), .B0(n4779), .B1(n3950), .Y(n4111) );
  OAI22XL U3890 ( .A0(n4756), .A1(n4024), .B0(n3949), .B1(n4112), .Y(n4110) );
  OAI22XL U3891 ( .A0(n4746), .A1(n3467), .B0(n2996), .B1(n4113), .Y(n4109) );
  OAI2BB2XL U3892 ( .B0(n2112), .B1(n4027), .A0N(N4278), .A1N(n4028), .Y(n4108) );
  OA22X1 U3893 ( .A0(n4029), .A1(n4813), .B0(n4114), .B1(n3440), .Y(n4104) );
  AOI222XL U3894 ( .A0(N2189), .A1(n4031), .B0(n4032), .B1(IM_Q[7]), .C0(N244), 
        .C1(n4018), .Y(n4114) );
  OA22X1 U3895 ( .A0(n4033), .A1(n4112), .B0(n4034), .B1(n4113), .Y(n4103) );
  CLKINVX1 U3896 ( .A(N3695), .Y(n4113) );
  CLKINVX1 U3897 ( .A(N3670), .Y(n4112) );
  OAI22XL U3898 ( .A0(n4746), .A1(n4035), .B0(n4779), .B1(n4036), .Y(n4102) );
  OR4X1 U3899 ( .A(n4115), .B(n4116), .C(n4117), .D(n4118), .Y(n1481) );
  OAI22XL U3900 ( .A0(n4812), .A1(n4029), .B0(n4119), .B1(n3440), .Y(n4118) );
  AOI222XL U3901 ( .A0(N2190), .A1(n4031), .B0(IM_Q[8]), .B1(n4032), .C0(N243), 
        .C1(n4018), .Y(n4119) );
  OAI21XL U3902 ( .A0(n4120), .A1(n3316), .B0(n4121), .Y(n4117) );
  AOI2BB2X1 U3903 ( .B0(n4018), .B1(N243), .A0N(n4122), .A1N(n3347), .Y(n4120)
         );
  NOR4X1 U3904 ( .A(n4123), .B(n4124), .C(n4125), .D(n4126), .Y(n4122) );
  OAI22XL U3905 ( .A0(n4812), .A1(n4023), .B0(n4778), .B1(n3950), .Y(n4126) );
  OAI22XL U3906 ( .A0(n4755), .A1(n4024), .B0(n3949), .B1(n4127), .Y(n4125) );
  OAI22XL U3907 ( .A0(n2083), .A1(n3467), .B0(n2996), .B1(n4128), .Y(n4124) );
  OAI2BB2XL U3908 ( .B0(n2111), .B1(n4027), .A0N(N4279), .A1N(n4028), .Y(n4123) );
  OAI22XL U3909 ( .A0(n4034), .A1(n4128), .B0(n4033), .B1(n4127), .Y(n4116) );
  CLKINVX1 U3910 ( .A(N3671), .Y(n4127) );
  CLKINVX1 U3911 ( .A(N3696), .Y(n4128) );
  OAI22XL U3912 ( .A0(n2083), .A1(n4035), .B0(n4778), .B1(n4036), .Y(n4115) );
  NAND4X1 U3913 ( .A(n4129), .B(n4130), .C(n4131), .D(n4132), .Y(n1480) );
  AOI221XL U3914 ( .A0(n4133), .A1(\IM_D_t[3][9] ), .B0(N2191), .B1(n4134), 
        .C0(n4016), .Y(n4132) );
  AOI222XL U3915 ( .A0(N242), .A1(n4135), .B0(N4280), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][9] ), .Y(n4131) );
  AOI222XL U3916 ( .A0(n4138), .A1(\IM_D_t[2][9] ), .B0(N3672), .B1(n4139), 
        .C0(N3697), .C1(n4140), .Y(n4130) );
  AOI222XL U3917 ( .A0(n4141), .A1(IM_Q[9]), .B0(n4142), .B1(n4977), .C0(n4143), .C1(\IM_D_t[0][9] ), .Y(n4129) );
  NAND4X1 U3918 ( .A(n4144), .B(n4145), .C(n4146), .D(n4147), .Y(n1479) );
  AOI221XL U3919 ( .A0(n4133), .A1(\IM_D_t[3][10] ), .B0(N2192), .B1(n4134), 
        .C0(n4016), .Y(n4147) );
  AOI222XL U3920 ( .A0(N241), .A1(n4135), .B0(N4281), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][10] ), .Y(n4146) );
  AOI222XL U3921 ( .A0(n4138), .A1(\IM_D_t[2][10] ), .B0(N3673), .B1(n4139), 
        .C0(N3698), .C1(n4140), .Y(n4145) );
  AOI222XL U3922 ( .A0(n4141), .A1(IM_Q[10]), .B0(n4142), .B1(n4976), .C0(
        n4143), .C1(\IM_D_t[0][10] ), .Y(n4144) );
  NAND4X1 U3923 ( .A(n4148), .B(n4149), .C(n4150), .D(n4151), .Y(n1478) );
  AOI221XL U3924 ( .A0(n4133), .A1(\IM_D_t[3][11] ), .B0(N2193), .B1(n4134), 
        .C0(n4016), .Y(n4151) );
  AOI222XL U3925 ( .A0(N240), .A1(n4135), .B0(N4282), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][11] ), .Y(n4150) );
  AOI222XL U3926 ( .A0(n4138), .A1(\IM_D_t[2][11] ), .B0(N3674), .B1(n4139), 
        .C0(N3699), .C1(n4140), .Y(n4149) );
  AOI222XL U3927 ( .A0(n4141), .A1(IM_Q[11]), .B0(n4142), .B1(n4975), .C0(
        n4143), .C1(\IM_D_t[0][11] ), .Y(n4148) );
  NAND4X1 U3928 ( .A(n4152), .B(n4153), .C(n4154), .D(n4155), .Y(n1477) );
  AOI221XL U3929 ( .A0(n4133), .A1(\IM_D_t[3][12] ), .B0(N2194), .B1(n4134), 
        .C0(n4016), .Y(n4155) );
  AOI222XL U3930 ( .A0(N239), .A1(n4135), .B0(N4283), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][12] ), .Y(n4154) );
  AOI222XL U3931 ( .A0(n4138), .A1(\IM_D_t[2][12] ), .B0(N3675), .B1(n4139), 
        .C0(N3700), .C1(n4140), .Y(n4153) );
  AOI222XL U3932 ( .A0(n4141), .A1(IM_Q[12]), .B0(n4142), .B1(n4974), .C0(
        n4143), .C1(\IM_D_t[0][12] ), .Y(n4152) );
  NAND4X1 U3933 ( .A(n4156), .B(n4157), .C(n4158), .D(n4159), .Y(n1476) );
  AOI221XL U3934 ( .A0(n4133), .A1(\IM_D_t[3][13] ), .B0(N2195), .B1(n4134), 
        .C0(n4016), .Y(n4159) );
  AOI222XL U3935 ( .A0(N238), .A1(n4135), .B0(N4284), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][13] ), .Y(n4158) );
  AOI222XL U3936 ( .A0(n4138), .A1(\IM_D_t[2][13] ), .B0(N3676), .B1(n4139), 
        .C0(N3701), .C1(n4140), .Y(n4157) );
  AOI222XL U3937 ( .A0(n4141), .A1(IM_Q[13]), .B0(n4142), .B1(n4973), .C0(
        n4143), .C1(\IM_D_t[0][13] ), .Y(n4156) );
  NAND4X1 U3938 ( .A(n4160), .B(n4161), .C(n4162), .D(n4163), .Y(n1475) );
  AOI221XL U3939 ( .A0(n4133), .A1(\IM_D_t[3][14] ), .B0(N2196), .B1(n4134), 
        .C0(n4016), .Y(n4163) );
  AOI222XL U3940 ( .A0(N237), .A1(n4135), .B0(N4285), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][14] ), .Y(n4162) );
  AOI222XL U3941 ( .A0(n4138), .A1(\IM_D_t[2][14] ), .B0(N3677), .B1(n4139), 
        .C0(N3702), .C1(n4140), .Y(n4161) );
  AOI222XL U3942 ( .A0(n4141), .A1(IM_Q[14]), .B0(n4142), .B1(n4972), .C0(
        n4143), .C1(\IM_D_t[0][14] ), .Y(n4160) );
  NAND4X1 U3943 ( .A(n4164), .B(n4165), .C(n4166), .D(n4167), .Y(n1474) );
  AOI221XL U3944 ( .A0(n4133), .A1(\IM_D_t[3][15] ), .B0(N2197), .B1(n4134), 
        .C0(n4016), .Y(n4167) );
  AOI222XL U3945 ( .A0(N236), .A1(n4135), .B0(N4286), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][15] ), .Y(n4166) );
  AOI222XL U3946 ( .A0(n4138), .A1(\IM_D_t[2][15] ), .B0(N3678), .B1(n4139), 
        .C0(N3703), .C1(n4140), .Y(n4165) );
  AOI222XL U3947 ( .A0(n4141), .A1(IM_Q[15]), .B0(n4142), .B1(n4971), .C0(
        n4143), .C1(\IM_D_t[0][15] ), .Y(n4164) );
  NAND4X1 U3948 ( .A(n4168), .B(n4169), .C(n4170), .D(n4171), .Y(n1473) );
  AOI221XL U3949 ( .A0(n4133), .A1(\IM_D_t[3][16] ), .B0(N2198), .B1(n4134), 
        .C0(n4016), .Y(n4171) );
  AOI222XL U3950 ( .A0(N235), .A1(n4135), .B0(N4287), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][16] ), .Y(n4170) );
  AOI222XL U3951 ( .A0(n4138), .A1(\IM_D_t[2][16] ), .B0(N3679), .B1(n4139), 
        .C0(N3704), .C1(n4140), .Y(n4169) );
  AOI222XL U3952 ( .A0(n4141), .A1(IM_Q[16]), .B0(n4142), .B1(n4970), .C0(
        n4143), .C1(\IM_D_t[0][16] ), .Y(n4168) );
  NAND4X1 U3953 ( .A(n4172), .B(n4173), .C(n4174), .D(n4175), .Y(n1472) );
  AOI221XL U3954 ( .A0(n4133), .A1(\IM_D_t[3][17] ), .B0(N2199), .B1(n4134), 
        .C0(n4016), .Y(n4175) );
  AOI222XL U3955 ( .A0(N234), .A1(n4135), .B0(N4288), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][17] ), .Y(n4174) );
  AOI222XL U3956 ( .A0(n4138), .A1(\IM_D_t[2][17] ), .B0(N3680), .B1(n4139), 
        .C0(N3705), .C1(n4140), .Y(n4173) );
  AOI222XL U3957 ( .A0(n4141), .A1(IM_Q[17]), .B0(n4142), .B1(n4969), .C0(
        n4143), .C1(\IM_D_t[0][17] ), .Y(n4172) );
  NAND4X1 U3958 ( .A(n4176), .B(n4177), .C(n4178), .D(n4179), .Y(n1471) );
  AOI221XL U3959 ( .A0(n4133), .A1(\IM_D_t[3][18] ), .B0(N2200), .B1(n4134), 
        .C0(n4016), .Y(n4179) );
  AOI222XL U3960 ( .A0(N233), .A1(n4135), .B0(N4289), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][18] ), .Y(n4178) );
  AOI222XL U3961 ( .A0(n4138), .A1(\IM_D_t[2][18] ), .B0(N3681), .B1(n4139), 
        .C0(N3706), .C1(n4140), .Y(n4177) );
  AOI222XL U3962 ( .A0(n4141), .A1(IM_Q[18]), .B0(n4142), .B1(n4968), .C0(
        n4143), .C1(\IM_D_t[0][18] ), .Y(n4176) );
  NAND4X1 U3963 ( .A(n4180), .B(n4181), .C(n4182), .D(n4183), .Y(n1470) );
  AOI221XL U3964 ( .A0(n4133), .A1(\IM_D_t[3][19] ), .B0(N2201), .B1(n4134), 
        .C0(n4016), .Y(n4183) );
  AOI222XL U3965 ( .A0(N232), .A1(n4135), .B0(N4290), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][19] ), .Y(n4182) );
  AOI222XL U3966 ( .A0(n4138), .A1(\IM_D_t[2][19] ), .B0(N3682), .B1(n4139), 
        .C0(N3707), .C1(n4140), .Y(n4181) );
  AOI222XL U3967 ( .A0(n4141), .A1(IM_Q[19]), .B0(n4142), .B1(n4967), .C0(
        n4143), .C1(\IM_D_t[0][19] ), .Y(n4180) );
  NAND4X1 U3968 ( .A(n4184), .B(n4185), .C(n4186), .D(n4187), .Y(n1469) );
  AOI221XL U3969 ( .A0(n4133), .A1(\IM_D_t[3][20] ), .B0(N2202), .B1(n4134), 
        .C0(n4016), .Y(n4187) );
  AOI222XL U3970 ( .A0(N231), .A1(n4135), .B0(N4291), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][20] ), .Y(n4186) );
  AOI222XL U3971 ( .A0(n4138), .A1(\IM_D_t[2][20] ), .B0(N3683), .B1(n4139), 
        .C0(N3708), .C1(n4140), .Y(n4185) );
  AOI222XL U3972 ( .A0(n4141), .A1(IM_Q[20]), .B0(n4142), .B1(n4966), .C0(
        n4143), .C1(\IM_D_t[0][20] ), .Y(n4184) );
  NAND4X1 U3973 ( .A(n4188), .B(n4189), .C(n4190), .D(n4191), .Y(n1468) );
  AOI221XL U3974 ( .A0(n4133), .A1(\IM_D_t[3][21] ), .B0(N2203), .B1(n4134), 
        .C0(n4016), .Y(n4191) );
  AOI222XL U3975 ( .A0(N230), .A1(n4135), .B0(N4292), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][21] ), .Y(n4190) );
  AOI222XL U3976 ( .A0(n4138), .A1(\IM_D_t[2][21] ), .B0(N3684), .B1(n4139), 
        .C0(N3709), .C1(n4140), .Y(n4189) );
  AOI222XL U3977 ( .A0(n4141), .A1(IM_Q[21]), .B0(n4142), .B1(n4965), .C0(
        n4143), .C1(\IM_D_t[0][21] ), .Y(n4188) );
  NAND4X1 U3978 ( .A(n4192), .B(n4193), .C(n4194), .D(n4195), .Y(n1467) );
  AOI221XL U3979 ( .A0(n4133), .A1(\IM_D_t[3][22] ), .B0(N2204), .B1(n4134), 
        .C0(n4016), .Y(n4195) );
  AOI222XL U3980 ( .A0(N229), .A1(n4135), .B0(N4293), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][22] ), .Y(n4194) );
  AOI222XL U3981 ( .A0(n4138), .A1(\IM_D_t[2][22] ), .B0(N3685), .B1(n4139), 
        .C0(N3710), .C1(n4140), .Y(n4193) );
  AOI222XL U3982 ( .A0(n4141), .A1(IM_Q[22]), .B0(n4142), .B1(n4964), .C0(
        n4143), .C1(\IM_D_t[0][22] ), .Y(n4192) );
  NAND4X1 U3983 ( .A(n4196), .B(n4197), .C(n4198), .D(n4199), .Y(n1466) );
  AOI221XL U3984 ( .A0(n4133), .A1(\IM_D_t[3][23] ), .B0(N2205), .B1(n4134), 
        .C0(n4016), .Y(n4199) );
  OAI22XL U3985 ( .A0(n3333), .A1(n3331), .B0(n3441), .B1(n3665), .Y(n4200) );
  AOI222XL U3986 ( .A0(N228), .A1(n4135), .B0(N4294), .B1(n4136), .C0(n4137), 
        .C1(\IM_D_t[1][23] ), .Y(n4198) );
  AOI222XL U3987 ( .A0(n4138), .A1(\IM_D_t[2][23] ), .B0(N3686), .B1(n4139), 
        .C0(N3711), .C1(n4140), .Y(n4197) );
  NAND2BX1 U3988 ( .AN(n3665), .B(n3441), .Y(n3477) );
  AOI211X1 U3989 ( .A0(n4205), .A1(n4209), .B0(n3645), .C0(n3446), .Y(n4208)
         );
  OAI22XL U3990 ( .A0(n3531), .A1(n3527), .B0(n3201), .B1(n3202), .Y(n3446) );
  OA21XL U3991 ( .A0(n4210), .A1(n3202), .B0(n4211), .Y(n4207) );
  NAND4BX1 U3992 ( .AN(n4212), .B(n4213), .C(n4214), .D(n4215), .Y(n1465) );
  AOI221XL U3993 ( .A0(N3164), .A1(n4014), .B0(n3410), .B1(n4216), .C0(n4016), 
        .Y(n4215) );
  MXI4X1 U3994 ( .A(n4219), .B(n4220), .C(n4221), .D(n4222), .S0(n4873), .S1(
        n4874), .Y(n4218) );
  AOI221XL U3995 ( .A0(CR_Q[11]), .A1(n4223), .B0(CR_Q[12]), .B1(n3787), .C0(
        n4224), .Y(n4222) );
  AO22X1 U3996 ( .A0(CR_Q[10]), .A1(n4225), .B0(CR_Q[9]), .B1(n3817), .Y(n4224) );
  AOI221XL U3997 ( .A0(CR_Q[3]), .A1(n4223), .B0(CR_Q[4]), .B1(n3787), .C0(
        n4226), .Y(n4221) );
  AO22X1 U3998 ( .A0(CR_Q[2]), .A1(n4225), .B0(CR_Q[1]), .B1(n3817), .Y(n4226)
         );
  AOI221XL U3999 ( .A0(CR_Q[7]), .A1(n4223), .B0(CR_Q[8]), .B1(n3787), .C0(
        n4227), .Y(n4220) );
  AO22X1 U4000 ( .A0(CR_Q[6]), .A1(n4225), .B0(CR_Q[5]), .B1(n3817), .Y(n4227)
         );
  NOR2X1 U4001 ( .A(n1424), .B(n4875), .Y(n3817) );
  CLKINVX1 U4002 ( .A(CR_Q[0]), .Y(n4219) );
  OAI2BB2XL U4003 ( .B0(n4228), .B1(n3347), .A0N(n4018), .A1N(N251), .Y(n4216)
         );
  NOR4X1 U4004 ( .A(n4229), .B(n4230), .C(n4231), .D(n4232), .Y(n4228) );
  OAI22XL U4005 ( .A0(n4834), .A1(n4023), .B0(n4786), .B1(n3950), .Y(n4232) );
  OAI22XL U4006 ( .A0(n4777), .A1(n4024), .B0(n3949), .B1(n4233), .Y(n4231) );
  OAI22XL U4007 ( .A0(n4753), .A1(n3467), .B0(n2996), .B1(n4234), .Y(n4230) );
  OAI2BB2XL U4008 ( .B0(n2133), .B1(n4027), .A0N(N4271), .A1N(n4028), .Y(n4229) );
  NOR2X1 U4009 ( .A(n4004), .B(n3306), .Y(n3373) );
  OA22X1 U4010 ( .A0(n4029), .A1(n4834), .B0(n4235), .B1(n3440), .Y(n4214) );
  AOI222XL U4011 ( .A0(N2182), .A1(n4031), .B0(IM_Q[0]), .B1(n4032), .C0(N251), 
        .C1(n4018), .Y(n4235) );
  NAND2X1 U4012 ( .A(n4236), .B(n3333), .Y(n3483) );
  CLKINVX1 U4013 ( .A(N2136), .Y(n3333) );
  NAND2X1 U4014 ( .A(N2136), .B(n4236), .Y(n3524) );
  CLKINVX1 U4015 ( .A(n4237), .Y(n3441) );
  AOI2BB1X1 U4016 ( .A0N(n4206), .A1N(n3316), .B0(n3645), .Y(n4240) );
  NAND2X1 U4017 ( .A(n3459), .B(n3458), .Y(n3645) );
  NOR3BXL U4018 ( .AN(n4241), .B(n4242), .C(n3646), .Y(n4206) );
  OAI21XL U4019 ( .A0(n4242), .A1(n3646), .B0(n3433), .Y(n4239) );
  CLKINVX1 U4020 ( .A(n3440), .Y(n3433) );
  CLKINVX1 U4021 ( .A(n4243), .Y(n3646) );
  CLKINVX1 U4022 ( .A(n3390), .Y(n4238) );
  OA22X1 U4023 ( .A0(n4033), .A1(n4233), .B0(n4034), .B1(n4234), .Y(n4213) );
  CLKINVX1 U4024 ( .A(N3688), .Y(n4234) );
  CLKINVX1 U4025 ( .A(N3663), .Y(n4233) );
  OAI22XL U4026 ( .A0(n4753), .A1(n4035), .B0(n4786), .B1(n4036), .Y(n4212) );
  OAI31XL U4027 ( .A0(n4237), .A1(n3440), .A2(n3442), .B0(n4204), .Y(n4244) );
  OAI21XL U4028 ( .A0(n3426), .A1(n3188), .B0(n3761), .Y(n4237) );
  NAND4X1 U4029 ( .A(n4245), .B(n4246), .C(n4247), .D(n4248), .Y(n1464) );
  AOI221XL U4030 ( .A0(n4249), .A1(IM_WEN), .B0(n4251), .B1(n3423), .C0(n4252), 
        .Y(n4248) );
  CLKINVX1 U4031 ( .A(n3476), .Y(n4252) );
  NAND4X1 U4032 ( .A(n3460), .B(n4211), .C(n4253), .D(n4254), .Y(n4249) );
  AOI211X1 U4033 ( .A0(n3360), .A1(n4255), .B0(n4256), .C0(n3210), .Y(n4254)
         );
  OAI31XL U4034 ( .A0(n3408), .A1(n3202), .A2(n3623), .B0(n3407), .Y(n4256) );
  NAND2X1 U4035 ( .A(n3449), .B(n3528), .Y(n3408) );
  OAI211X1 U4036 ( .A0(n3347), .A1(n4023), .B0(n4241), .C0(n4210), .Y(n4255)
         );
  NOR3X1 U4037 ( .A(n3390), .B(n3423), .C(n3370), .Y(n4253) );
  NOR2X1 U4038 ( .A(n3798), .B(n3531), .Y(n3390) );
  CLKINVX1 U4039 ( .A(n3391), .Y(n3460) );
  NOR2X1 U4040 ( .A(n4243), .B(n3384), .Y(n3391) );
  NOR2X1 U4041 ( .A(n3360), .B(n3319), .Y(n3384) );
  NOR2BX1 U4042 ( .AN(n3289), .B(n3413), .Y(n4247) );
  NOR2X1 U4043 ( .A(n3647), .B(n3457), .Y(n3413) );
  NAND4X1 U4044 ( .A(n4223), .B(n4258), .C(N6484), .D(count[3]), .Y(n3647) );
  OAI31XL U4045 ( .A0(n4259), .A1(n3372), .A2(IM_WEN), .B0(n3371), .Y(n4246)
         );
  OAI31XL U4046 ( .A0(n4259), .A1(n3236), .A2(n3235), .B0(n3210), .Y(n4245) );
  NAND4X1 U4047 ( .A(n3259), .B(n4260), .C(n3258), .D(n4261), .Y(n4259) );
  NOR3X1 U4048 ( .A(n3239), .B(n3238), .C(n3237), .Y(n4261) );
  MXI2X1 U4049 ( .A(n4717), .B(n3806), .S0(n4262), .Y(n1463) );
  MXI2X1 U4050 ( .A(n4718), .B(n3808), .S0(n4262), .Y(n1462) );
  MXI2X1 U4051 ( .A(n4719), .B(n3809), .S0(n4262), .Y(n1461) );
  MXI2X1 U4052 ( .A(n4720), .B(n3810), .S0(n4262), .Y(n1460) );
  MXI2X1 U4053 ( .A(n4721), .B(n3811), .S0(n4262), .Y(n1459) );
  CLKINVX1 U4054 ( .A(IM_Q[15]), .Y(n3811) );
  MXI2X1 U4055 ( .A(n4722), .B(n3812), .S0(n4262), .Y(n1458) );
  MXI2X1 U4056 ( .A(n4723), .B(n3813), .S0(n4262), .Y(n1457) );
  CLKINVX1 U4057 ( .A(IM_Q[13]), .Y(n3813) );
  MXI2X1 U4058 ( .A(n4724), .B(n3814), .S0(n4262), .Y(n1456) );
  MXI2X1 U4059 ( .A(n4725), .B(n3815), .S0(n4262), .Y(n1455) );
  MXI2X1 U4060 ( .A(n4726), .B(n3816), .S0(n4262), .Y(n1454) );
  MXI2X1 U4061 ( .A(n4710), .B(n3299), .S0(n4262), .Y(n1451) );
  CLKINVX1 U4062 ( .A(IM_Q[7]), .Y(n3299) );
  MXI2X1 U4063 ( .A(n4711), .B(n3779), .S0(n4262), .Y(n1450) );
  CLKINVX1 U4064 ( .A(IM_Q[6]), .Y(n3779) );
  CLKINVX1 U4065 ( .A(IM_Q[5]), .Y(n3771) );
  CLKINVX1 U4066 ( .A(IM_Q[4]), .Y(n3773) );
  CLKINVX1 U4067 ( .A(IM_Q[3]), .Y(n3775) );
  NOR2X1 U4068 ( .A(n3354), .B(n3357), .Y(n3476) );
  CLKINVX1 U4069 ( .A(n3406), .Y(n3369) );
  NOR4X1 U4070 ( .A(n4269), .B(n4270), .C(n4271), .D(n4272), .Y(n4268) );
  AO22X1 U4071 ( .A0(n3210), .A1(n4273), .B0(n3371), .B1(n4274), .Y(n4272) );
  AOI222XL U4072 ( .A0(N647), .A1(n3237), .B0(N511), .B1(n3254), .C0(N551), 
        .C1(n3257), .Y(n4277) );
  OAI211X1 U4073 ( .A0(n3270), .A1(n4278), .B0(n4279), .C0(n4280), .Y(n4273)
         );
  AOI222XL U4074 ( .A0(N1359), .A1(n3237), .B0(N1282), .B1(n3235), .C0(N490), 
        .C1(n3236), .Y(n4280) );
  NAND2X1 U4075 ( .A(N1444), .B(n3238), .Y(n4279) );
  OAI22XL U4076 ( .A0(n3694), .A1(n3248), .B0(n3615), .B1(n3246), .Y(n4271) );
  AOI221XL U4077 ( .A0(N2788), .A1(n3560), .B0(N2853), .B1(n3561), .C0(n4281), 
        .Y(n3615) );
  MXI2X1 U4078 ( .A(N3735), .B(N2321), .S0(n3069), .Y(n3694) );
  AO22X1 U4079 ( .A0(count[3]), .A1(n3354), .B0(N3735), .B1(n3195), .Y(n4270)
         );
  OAI222XL U4080 ( .A0(n3284), .A1(n4275), .B0(n4282), .B1(n2983), .C0(n3286), 
        .C1(n4278), .Y(n4269) );
  CLKINVX1 U4081 ( .A(N947), .Y(n4278) );
  CLKINVX1 U4082 ( .A(N810), .Y(n4275) );
  AOI211X1 U4083 ( .A0(n3212), .A1(n4283), .B0(n4284), .C0(n4285), .Y(n4267)
         );
  OAI22XL U4084 ( .A0(n3574), .A1(n3295), .B0(n3741), .B1(n3297), .Y(n4285) );
  MXI2X1 U4085 ( .A(N2321), .B(N3735), .S0(n3069), .Y(n3741) );
  AOI221XL U4086 ( .A0(N4979), .A1(n3560), .B0(N5024), .B1(n3561), .C0(n4281), 
        .Y(n3574) );
  NOR2X1 U4087 ( .A(n3623), .B(n4841), .Y(n4281) );
  AO22X1 U4088 ( .A0(n4286), .A1(N490), .B0(N870), .B1(n3291), .Y(n4284) );
  NAND4X1 U4089 ( .A(n4287), .B(n4288), .C(n4289), .D(n4290), .Y(n4283) );
  AOI222XL U4090 ( .A0(N3755), .A1(n3218), .B0(n3219), .B1(IM_A[3]), .C0(N3620), .C1(n3220), .Y(n4290) );
  AOI22X1 U4091 ( .A0(N3735), .A1(n3221), .B0(N3735), .B1(n3222), .Y(n4289) );
  AOI22X1 U4092 ( .A0(N4457), .A1(n3223), .B0(N4179), .B1(n3224), .Y(n4288) );
  AOI22X1 U4093 ( .A0(N1027), .A1(n3292), .B0(n3243), .B1(N2321), .Y(n4266) );
  AOI2BB2X1 U4094 ( .B0(N6553), .B1(n3240), .A0N(n3290), .A1N(n4841), .Y(n4265) );
  NAND4BX1 U4095 ( .AN(n4292), .B(n4293), .C(n4294), .D(n4295), .Y(n1442) );
  AND4X1 U4096 ( .A(n4296), .B(n4297), .C(n4298), .D(n4299), .Y(n4295) );
  AOI222XL U4097 ( .A0(N512), .A1(n4300), .B0(n3354), .B1(count[4]), .C0(n3195), .C1(N3736), .Y(n4299) );
  AOI222XL U4098 ( .A0(N1360), .A1(n4301), .B0(N552), .B1(n4302), .C0(N1283), 
        .C1(n4303), .Y(n4298) );
  AOI222XL U4099 ( .A0(N713), .A1(n4304), .B0(N648), .B1(n3013), .C0(N1445), 
        .C1(n4306), .Y(n4297) );
  OA22X1 U4100 ( .A0(n3248), .A1(n3685), .B0(n3626), .B1(n3246), .Y(n4296) );
  AOI221XL U4101 ( .A0(N2789), .A1(n3560), .B0(N2854), .B1(n3561), .C0(n4307), 
        .Y(n3626) );
  MXI2X1 U4102 ( .A(N3736), .B(N2322), .S0(n3069), .Y(n3685) );
  AOI2BB2X1 U4103 ( .B0(N6554), .B1(n3240), .A0N(n3290), .A1N(n4840), .Y(n4294) );
  AOI222XL U4104 ( .A0(n3243), .A1(N2322), .B0(N1028), .B1(n3292), .C0(N948), 
        .C1(n4308), .Y(n4293) );
  OAI211X1 U4105 ( .A0(n4309), .A1(n3436), .B0(n4310), .C0(n4311), .Y(n4292)
         );
  AOI222XL U4106 ( .A0(N871), .A1(n3291), .B0(n3208), .B1(n3563), .C0(n3241), 
        .C1(n3732), .Y(n4311) );
  CLKMX2X2 U4107 ( .A(N3736), .B(N2322), .S0(n3381), .Y(n3732) );
  CLKINVX1 U4108 ( .A(n4312), .Y(n3563) );
  AOI221XL U4109 ( .A0(N4980), .A1(n3560), .B0(N5025), .B1(n3561), .C0(n4307), 
        .Y(n4312) );
  NOR2X1 U4110 ( .A(n3623), .B(n4840), .Y(n4307) );
  AOI22X1 U4111 ( .A0(N811), .A1(n4313), .B0(N491), .B1(n4314), .Y(n4310) );
  AND4X1 U4112 ( .A(n4315), .B(n4316), .C(n4317), .D(n4318), .Y(n4309) );
  AOI222XL U4113 ( .A0(N3756), .A1(n3218), .B0(n3219), .B1(IM_A[4]), .C0(N3621), .C1(n3220), .Y(n4318) );
  AOI22X1 U4114 ( .A0(N3736), .A1(n3221), .B0(N3736), .B1(n3222), .Y(n4317) );
  AOI22X1 U4115 ( .A0(N4458), .A1(n3223), .B0(N4180), .B1(n3224), .Y(n4316) );
  AOI22X1 U4116 ( .A0(N4110), .A1(n2998), .B0(N4368), .B1(n3226), .Y(n4315) );
  NAND4BX1 U4117 ( .AN(n4320), .B(n4321), .C(n4322), .D(n4323), .Y(n1441) );
  AND4X1 U4118 ( .A(n4324), .B(n4325), .C(n4326), .D(n4327), .Y(n4323) );
  AOI222XL U4119 ( .A0(N513), .A1(n4300), .B0(n3354), .B1(n3424), .C0(n3195), 
        .C1(N3737), .Y(n4327) );
  AOI222XL U4120 ( .A0(N1361), .A1(n4301), .B0(N553), .B1(n4302), .C0(N1284), 
        .C1(n4303), .Y(n4326) );
  AOI222XL U4121 ( .A0(N714), .A1(n4304), .B0(N649), .B1(n3013), .C0(N1446), 
        .C1(n4306), .Y(n4325) );
  OA22X1 U4122 ( .A0(n3248), .A1(n3679), .B0(n3636), .B1(n3246), .Y(n4324) );
  AOI221XL U4123 ( .A0(N2790), .A1(n3560), .B0(N2855), .B1(n3561), .C0(n4328), 
        .Y(n3636) );
  AOI2BB2X1 U4124 ( .B0(N6555), .B1(n3240), .A0N(n3290), .A1N(n4839), .Y(n4322) );
  AOI222XL U4125 ( .A0(n3243), .A1(N2323), .B0(N1029), .B1(n3292), .C0(N949), 
        .C1(n4308), .Y(n4321) );
  OAI211X1 U4126 ( .A0(n4329), .A1(n3436), .B0(n4330), .C0(n4331), .Y(n4320)
         );
  AOI222XL U4127 ( .A0(N872), .A1(n3291), .B0(n3208), .B1(n4332), .C0(n3241), 
        .C1(n3726), .Y(n4331) );
  CLKMX2X2 U4128 ( .A(N3737), .B(N2323), .S0(n3381), .Y(n3726) );
  CLKINVX1 U4129 ( .A(n3554), .Y(n4332) );
  AOI221XL U4130 ( .A0(N4981), .A1(n3560), .B0(N5026), .B1(n3561), .C0(n4328), 
        .Y(n3554) );
  NOR2X1 U4131 ( .A(n3623), .B(n4839), .Y(n4328) );
  AOI22X1 U4132 ( .A0(N812), .A1(n4313), .B0(N492), .B1(n4314), .Y(n4330) );
  AND4X1 U4133 ( .A(n4333), .B(n4334), .C(n4335), .D(n4336), .Y(n4329) );
  AOI222XL U4134 ( .A0(N3757), .A1(n3218), .B0(n3219), .B1(IM_A[5]), .C0(N3622), .C1(n3220), .Y(n4336) );
  AOI22X1 U4135 ( .A0(N3737), .A1(n3221), .B0(N3737), .B1(n3222), .Y(n4335) );
  AOI22X1 U4136 ( .A0(N4459), .A1(n3223), .B0(N4181), .B1(n3224), .Y(n4334) );
  AOI22X1 U4137 ( .A0(N4111), .A1(n2998), .B0(N4369), .B1(n3226), .Y(n4333) );
  NAND4BX1 U4138 ( .AN(n4338), .B(n4339), .C(n4340), .D(n4341), .Y(n1440) );
  AND4X1 U4139 ( .A(n4342), .B(n4343), .C(n4344), .D(n4345), .Y(n4341) );
  AOI222XL U4140 ( .A0(N514), .A1(n4300), .B0(n3354), .B1(n3425), .C0(n3195), 
        .C1(N3738), .Y(n4345) );
  AOI222XL U4141 ( .A0(N1362), .A1(n4301), .B0(N554), .B1(n4302), .C0(N1285), 
        .C1(n4303), .Y(n4344) );
  AOI222XL U4142 ( .A0(N715), .A1(n4304), .B0(N650), .B1(n3013), .C0(N1447), 
        .C1(n4306), .Y(n4343) );
  OA22X1 U4143 ( .A0(n3248), .A1(n3688), .B0(n3627), .B1(n3246), .Y(n4342) );
  AOI221XL U4144 ( .A0(N2791), .A1(n3560), .B0(N2856), .B1(n3561), .C0(n4346), 
        .Y(n3627) );
  AOI2BB2X1 U4145 ( .B0(N6556), .B1(n3240), .A0N(n3290), .A1N(n4838), .Y(n4340) );
  AOI222XL U4146 ( .A0(n3243), .A1(N2324), .B0(N1030), .B1(n3292), .C0(N950), 
        .C1(n4308), .Y(n4339) );
  OAI211X1 U4147 ( .A0(n4347), .A1(n3436), .B0(n4348), .C0(n4349), .Y(n4338)
         );
  AOI222XL U4148 ( .A0(N873), .A1(n3291), .B0(n3208), .B1(n4350), .C0(n3241), 
        .C1(n3735), .Y(n4349) );
  CLKMX2X2 U4149 ( .A(N3738), .B(N2324), .S0(n3381), .Y(n3735) );
  CLKINVX1 U4150 ( .A(n3568), .Y(n4350) );
  AOI221XL U4151 ( .A0(N4982), .A1(n3560), .B0(N5027), .B1(n3561), .C0(n4346), 
        .Y(n3568) );
  NOR2X1 U4152 ( .A(n3623), .B(n4838), .Y(n4346) );
  AOI22X1 U4153 ( .A0(N813), .A1(n4313), .B0(N493), .B1(n4314), .Y(n4348) );
  AND4X1 U4154 ( .A(n4351), .B(n4352), .C(n4353), .D(n4354), .Y(n4347) );
  AOI222XL U4155 ( .A0(N3758), .A1(n3218), .B0(n3219), .B1(IM_A[6]), .C0(N3623), .C1(n3220), .Y(n4354) );
  AOI22X1 U4156 ( .A0(N3738), .A1(n3221), .B0(N3738), .B1(n3222), .Y(n4353) );
  AOI22X1 U4157 ( .A0(N4112), .A1(n2998), .B0(N4370), .B1(n3226), .Y(n4351) );
  NAND4BX1 U4158 ( .AN(n4356), .B(n4357), .C(n4358), .D(n4359), .Y(n1439) );
  AND4X1 U4159 ( .A(n4360), .B(n4361), .C(n4362), .D(n4363), .Y(n4359) );
  AOI222XL U4160 ( .A0(N515), .A1(n4300), .B0(n3354), .B1(n3426), .C0(n3195), 
        .C1(N3739), .Y(n4363) );
  AOI222XL U4161 ( .A0(N1363), .A1(n4301), .B0(N555), .B1(n4302), .C0(N1286), 
        .C1(n4303), .Y(n4362) );
  AOI222XL U4162 ( .A0(N716), .A1(n4304), .B0(N651), .B1(n3013), .C0(N1448), 
        .C1(n4306), .Y(n4361) );
  OA22X1 U4163 ( .A0(n3248), .A1(n3689), .B0(n3628), .B1(n3246), .Y(n4360) );
  AOI221XL U4164 ( .A0(N2792), .A1(n3560), .B0(N2857), .B1(n3561), .C0(n4364), 
        .Y(n3628) );
  MXI2X1 U4165 ( .A(N3739), .B(N2325), .S0(n3069), .Y(n3689) );
  AOI2BB2X1 U4166 ( .B0(N6557), .B1(n3240), .A0N(n3290), .A1N(n4837), .Y(n4358) );
  AOI222XL U4167 ( .A0(n3243), .A1(N2325), .B0(N1031), .B1(n3292), .C0(N951), 
        .C1(n4308), .Y(n4357) );
  OAI211X1 U4168 ( .A0(n4365), .A1(n3436), .B0(n4366), .C0(n4367), .Y(n4356)
         );
  AOI222XL U4169 ( .A0(N874), .A1(n3291), .B0(n3208), .B1(n4368), .C0(n3241), 
        .C1(n3736), .Y(n4367) );
  CLKMX2X2 U4170 ( .A(N3739), .B(N2325), .S0(n3381), .Y(n3736) );
  CLKINVX1 U4171 ( .A(n3569), .Y(n4368) );
  AOI221XL U4172 ( .A0(N4983), .A1(n3560), .B0(N5028), .B1(n3561), .C0(n4364), 
        .Y(n3569) );
  NOR2X1 U4173 ( .A(n3623), .B(n4837), .Y(n4364) );
  AOI22X1 U4174 ( .A0(N814), .A1(n4313), .B0(N494), .B1(n4314), .Y(n4366) );
  AND4X1 U4175 ( .A(n4369), .B(n4370), .C(n4371), .D(n4372), .Y(n4365) );
  AOI222XL U4176 ( .A0(N3759), .A1(n3218), .B0(n3219), .B1(IM_A[7]), .C0(N3624), .C1(n3220), .Y(n4372) );
  AOI22X1 U4177 ( .A0(N3739), .A1(n3221), .B0(N3739), .B1(n3222), .Y(n4371) );
  NAND4BX1 U4178 ( .AN(n4374), .B(n4375), .C(n4376), .D(n4377), .Y(n1438) );
  AOI222XL U4179 ( .A0(N6558), .A1(n3240), .B0(N815), .B1(n3001), .C0(n3243), 
        .C1(N2326), .Y(n4377) );
  NOR3BXL U4180 ( .AN(n4378), .B(n4379), .C(n4380), .Y(n4376) );
  OAI22XL U4181 ( .A0(n4836), .A1(n4381), .B0(n4382), .B1(n4383), .Y(n4380) );
  CLKINVX1 U4182 ( .A(N3740), .Y(n4383) );
  OAI22XL U4183 ( .A0(n3705), .A1(n3248), .B0(n3604), .B1(n3246), .Y(n4379) );
  AOI221XL U4184 ( .A0(N2793), .A1(n3560), .B0(N2858), .B1(n3561), .C0(n4384), 
        .Y(n3604) );
  MXI2X1 U4185 ( .A(N3740), .B(N2326), .S0(n3069), .Y(n3705) );
  AOI222XL U4186 ( .A0(n3208), .A1(n3585), .B0(N495), .B1(n4314), .C0(n3241), 
        .C1(n3752), .Y(n4378) );
  CLKMX2X2 U4187 ( .A(N3740), .B(N2326), .S0(n3381), .Y(n3752) );
  CLKINVX1 U4188 ( .A(n4385), .Y(n3585) );
  AOI221XL U4189 ( .A0(N4984), .A1(n3560), .B0(N5029), .B1(n3561), .C0(n4384), 
        .Y(n4385) );
  NOR2X1 U4190 ( .A(n3623), .B(n4836), .Y(n4384) );
  AOI222XL U4191 ( .A0(N952), .A1(n4308), .B0(N875), .B1(n3291), .C0(N1032), 
        .C1(n3292), .Y(n4375) );
  NAND4X1 U4192 ( .A(n4386), .B(n4387), .C(n4388), .D(n4389), .Y(n4374) );
  AND3X1 U4193 ( .A(n4390), .B(n4391), .C(n4392), .Y(n4389) );
  AOI222XL U4194 ( .A0(N717), .A1(n4304), .B0(N652), .B1(n3013), .C0(N1449), 
        .C1(n4306), .Y(n4392) );
  AOI22X1 U4195 ( .A0(N516), .A1(n4300), .B0(N556), .B1(n4302), .Y(n4391) );
  AOI22X1 U4196 ( .A0(N1287), .A1(n4303), .B0(N1364), .B1(n4301), .Y(n4390) );
  AOI222XL U4197 ( .A0(N4372), .A1(n4393), .B0(N4184), .B1(n4394), .C0(N4114), 
        .C1(n3000), .Y(n4388) );
  NAND4BX1 U4198 ( .AN(n4400), .B(n4401), .C(n4402), .D(n4403), .Y(n1437) );
  AOI222XL U4199 ( .A0(N6559), .A1(n3240), .B0(N816), .B1(n3001), .C0(n3243), 
        .C1(N2327), .Y(n4403) );
  NOR3BXL U4200 ( .AN(n4404), .B(n4405), .C(n4406), .Y(n4402) );
  OAI22XL U4201 ( .A0(n4835), .A1(n4381), .B0(n4382), .B1(N3741), .Y(n4406) );
  OAI22XL U4202 ( .A0(n3707), .A1(n3248), .B0(n3601), .B1(n3246), .Y(n4405) );
  AOI221XL U4203 ( .A0(N2794), .A1(n3560), .B0(N2859), .B1(n3561), .C0(n4407), 
        .Y(n3601) );
  MXI2X1 U4204 ( .A(N2413), .B(N2327), .S0(n3069), .Y(n3707) );
  AOI222XL U4205 ( .A0(n3208), .A1(n3587), .B0(N496), .B1(n4314), .C0(n3241), 
        .C1(n3754), .Y(n4404) );
  CLKMX2X2 U4206 ( .A(N2413), .B(N2327), .S0(n3381), .Y(n3754) );
  CLKINVX1 U4207 ( .A(n4408), .Y(n3587) );
  AOI221XL U4208 ( .A0(N4985), .A1(n3560), .B0(N5030), .B1(n3561), .C0(n4407), 
        .Y(n4408) );
  NOR2X1 U4209 ( .A(n3623), .B(n4835), .Y(n4407) );
  AOI222XL U4210 ( .A0(N953), .A1(n4308), .B0(N876), .B1(n3291), .C0(N1033), 
        .C1(n3292), .Y(n4401) );
  NAND4X1 U4211 ( .A(n4409), .B(n4410), .C(n4411), .D(n4412), .Y(n4400) );
  AND3X1 U4212 ( .A(n4413), .B(n4414), .C(n4415), .Y(n4412) );
  AOI222XL U4213 ( .A0(N718), .A1(n4304), .B0(N653), .B1(n3013), .C0(N1450), 
        .C1(n4306), .Y(n4415) );
  AOI22X1 U4214 ( .A0(N517), .A1(n4300), .B0(N557), .B1(n4302), .Y(n4414) );
  AOI22X1 U4215 ( .A0(N1288), .A1(n4303), .B0(N1365), .B1(n4301), .Y(n4413) );
  AOI222XL U4216 ( .A0(N4373), .A1(n4393), .B0(N4185), .B1(n4394), .C0(N4115), 
        .C1(n3000), .Y(n4411) );
  NAND4BX1 U4217 ( .AN(n4416), .B(n4417), .C(n4418), .D(n4419), .Y(n1436) );
  AOI222XL U4218 ( .A0(N6560), .A1(n3240), .B0(N817), .B1(n3001), .C0(n3243), 
        .C1(N2328), .Y(n4419) );
  NOR3BXL U4219 ( .AN(n4420), .B(n4421), .C(n4422), .Y(n4418) );
  OAI22XL U4220 ( .A0(n4853), .A1(n4381), .B0(n4382), .B1(n4423), .Y(n4422) );
  CLKINVX1 U4221 ( .A(N2414), .Y(n4423) );
  OAI22XL U4222 ( .A0(n3706), .A1(n3248), .B0(n3605), .B1(n3246), .Y(n4421) );
  AOI221XL U4223 ( .A0(N2795), .A1(n3560), .B0(N2860), .B1(n3561), .C0(n4424), 
        .Y(n3605) );
  MXI2X1 U4224 ( .A(N2414), .B(N2328), .S0(n3069), .Y(n3706) );
  AOI222XL U4225 ( .A0(n3208), .A1(n3586), .B0(N497), .B1(n4314), .C0(n3241), 
        .C1(n3753), .Y(n4420) );
  CLKMX2X2 U4226 ( .A(N2414), .B(N2328), .S0(n3381), .Y(n3753) );
  CLKINVX1 U4227 ( .A(n4425), .Y(n3586) );
  AOI221XL U4228 ( .A0(N4986), .A1(n3560), .B0(N5031), .B1(n3561), .C0(n4424), 
        .Y(n4425) );
  NOR2X1 U4229 ( .A(n3623), .B(n4853), .Y(n4424) );
  AOI222XL U4230 ( .A0(N954), .A1(n4308), .B0(N877), .B1(n3291), .C0(N1034), 
        .C1(n3292), .Y(n4417) );
  NAND4X1 U4231 ( .A(n4426), .B(n4427), .C(n4428), .D(n4429), .Y(n4416) );
  AND3X1 U4232 ( .A(n4430), .B(n4431), .C(n4432), .Y(n4429) );
  AOI222XL U4233 ( .A0(N719), .A1(n4304), .B0(N654), .B1(n3013), .C0(N1451), 
        .C1(n4306), .Y(n4432) );
  AOI22X1 U4234 ( .A0(N518), .A1(n4300), .B0(N558), .B1(n4302), .Y(n4431) );
  AOI22X1 U4235 ( .A0(N1289), .A1(n4303), .B0(N1366), .B1(n4301), .Y(n4430) );
  AOI222XL U4236 ( .A0(N4374), .A1(n4393), .B0(N4186), .B1(n4394), .C0(N4116), 
        .C1(n3000), .Y(n4428) );
  NAND4BX1 U4237 ( .AN(n4433), .B(n4434), .C(n4435), .D(n4436), .Y(n1435) );
  AOI222XL U4238 ( .A0(N6561), .A1(n3240), .B0(N818), .B1(n3001), .C0(n3243), 
        .C1(N2329), .Y(n4436) );
  NOR3BXL U4239 ( .AN(n4437), .B(n4438), .C(n4439), .Y(n4435) );
  OAI22XL U4240 ( .A0(n4852), .A1(n4381), .B0(n4382), .B1(n4440), .Y(n4439) );
  CLKINVX1 U4241 ( .A(N2415), .Y(n4440) );
  OAI22XL U4242 ( .A0(n3710), .A1(n3248), .B0(n3606), .B1(n3246), .Y(n4438) );
  AOI221XL U4243 ( .A0(N2796), .A1(n3560), .B0(N2861), .B1(n3561), .C0(n4441), 
        .Y(n3606) );
  MXI2X1 U4244 ( .A(N2415), .B(N2329), .S0(n3069), .Y(n3710) );
  AOI222XL U4245 ( .A0(n3208), .A1(n4442), .B0(N498), .B1(n4314), .C0(n3241), 
        .C1(n3757), .Y(n4437) );
  CLKMX2X2 U4246 ( .A(N2415), .B(N2329), .S0(n3381), .Y(n3757) );
  CLKINVX1 U4247 ( .A(n3590), .Y(n4442) );
  AOI221XL U4248 ( .A0(N4987), .A1(n3560), .B0(N5032), .B1(n3561), .C0(n4441), 
        .Y(n3590) );
  NOR2X1 U4249 ( .A(n3623), .B(n4852), .Y(n4441) );
  AOI222XL U4250 ( .A0(N955), .A1(n4308), .B0(N878), .B1(n3291), .C0(N1035), 
        .C1(n3292), .Y(n4434) );
  NAND4X1 U4251 ( .A(n4443), .B(n4444), .C(n4445), .D(n4446), .Y(n4433) );
  AND3X1 U4252 ( .A(n4447), .B(n4448), .C(n4449), .Y(n4446) );
  AOI222XL U4253 ( .A0(N720), .A1(n4304), .B0(N655), .B1(n3013), .C0(N1452), 
        .C1(n4306), .Y(n4449) );
  AOI22X1 U4254 ( .A0(N519), .A1(n4300), .B0(N559), .B1(n4302), .Y(n4448) );
  AOI22X1 U4255 ( .A0(N1290), .A1(n4303), .B0(N1367), .B1(n4301), .Y(n4447) );
  AOI222XL U4256 ( .A0(N4375), .A1(n4393), .B0(N4187), .B1(n4394), .C0(N4117), 
        .C1(n3000), .Y(n4445) );
  NAND4BX1 U4257 ( .AN(n4450), .B(n4451), .C(n4452), .D(n4453), .Y(n1434) );
  AOI222XL U4258 ( .A0(N6562), .A1(n3240), .B0(N819), .B1(n3001), .C0(n3243), 
        .C1(N2330), .Y(n4453) );
  NOR3BXL U4259 ( .AN(n4454), .B(n4455), .C(n4456), .Y(n4452) );
  OAI22XL U4260 ( .A0(n4851), .A1(n4381), .B0(n4382), .B1(n4457), .Y(n4456) );
  CLKINVX1 U4261 ( .A(N2416), .Y(n4457) );
  OAI22XL U4262 ( .A0(n3696), .A1(n3248), .B0(n3612), .B1(n3246), .Y(n4455) );
  AOI221XL U4263 ( .A0(N2797), .A1(n3560), .B0(N2862), .B1(n3561), .C0(n4458), 
        .Y(n3612) );
  MXI2X1 U4264 ( .A(N2416), .B(N2330), .S0(n3069), .Y(n3696) );
  AOI222XL U4265 ( .A0(n3208), .A1(n3576), .B0(N499), .B1(n4314), .C0(n3241), 
        .C1(n3743), .Y(n4454) );
  CLKMX2X2 U4266 ( .A(N2416), .B(N2330), .S0(n3381), .Y(n3743) );
  CLKINVX1 U4267 ( .A(n4459), .Y(n3576) );
  AOI221XL U4268 ( .A0(N4988), .A1(n3560), .B0(N5033), .B1(n3561), .C0(n4458), 
        .Y(n4459) );
  NOR2X1 U4269 ( .A(n3623), .B(n4851), .Y(n4458) );
  AOI222XL U4270 ( .A0(N956), .A1(n4308), .B0(N879), .B1(n3291), .C0(N1036), 
        .C1(n3292), .Y(n4451) );
  NAND4X1 U4271 ( .A(n4460), .B(n4461), .C(n4462), .D(n4463), .Y(n4450) );
  AND3X1 U4272 ( .A(n4464), .B(n4465), .C(n4466), .Y(n4463) );
  AOI222XL U4273 ( .A0(N721), .A1(n4304), .B0(N656), .B1(n3013), .C0(N1453), 
        .C1(n4306), .Y(n4466) );
  AOI22X1 U4274 ( .A0(N520), .A1(n4300), .B0(N560), .B1(n4302), .Y(n4465) );
  AOI22X1 U4275 ( .A0(N1291), .A1(n4303), .B0(N1368), .B1(n4301), .Y(n4464) );
  AOI222XL U4276 ( .A0(N4376), .A1(n4393), .B0(N4188), .B1(n4394), .C0(N4118), 
        .C1(n3000), .Y(n4462) );
  NAND4BX1 U4277 ( .AN(n4467), .B(n4468), .C(n4469), .D(n4470), .Y(n1433) );
  AOI222XL U4278 ( .A0(N6563), .A1(n3240), .B0(N820), .B1(n3001), .C0(n3243), 
        .C1(N2331), .Y(n4470) );
  NOR3BXL U4279 ( .AN(n4471), .B(n4472), .C(n4473), .Y(n4469) );
  OAI22XL U4280 ( .A0(n4850), .A1(n4381), .B0(n4382), .B1(n4474), .Y(n4473) );
  CLKINVX1 U4281 ( .A(N2417), .Y(n4474) );
  OAI22XL U4282 ( .A0(n3695), .A1(n3248), .B0(n3616), .B1(n3246), .Y(n4472) );
  AOI221XL U4283 ( .A0(N2798), .A1(n3560), .B0(N2863), .B1(n3561), .C0(n4475), 
        .Y(n3616) );
  MXI2X1 U4284 ( .A(N2417), .B(N2331), .S0(n3069), .Y(n3695) );
  AOI222XL U4285 ( .A0(n3208), .A1(n3575), .B0(N500), .B1(n4314), .C0(n3241), 
        .C1(n3742), .Y(n4471) );
  CLKMX2X2 U4286 ( .A(N2417), .B(N2331), .S0(n3381), .Y(n3742) );
  CLKINVX1 U4287 ( .A(n4476), .Y(n3575) );
  AOI221XL U4288 ( .A0(N4989), .A1(n3560), .B0(N5034), .B1(n3561), .C0(n4475), 
        .Y(n4476) );
  NOR2X1 U4289 ( .A(n3623), .B(n4850), .Y(n4475) );
  AOI222XL U4290 ( .A0(N957), .A1(n4308), .B0(N880), .B1(n3291), .C0(N1037), 
        .C1(n3292), .Y(n4468) );
  NAND4X1 U4291 ( .A(n4477), .B(n4478), .C(n4479), .D(n4480), .Y(n4467) );
  AND3X1 U4292 ( .A(n4481), .B(n4482), .C(n4483), .Y(n4480) );
  AOI222XL U4293 ( .A0(N722), .A1(n4304), .B0(N657), .B1(n3013), .C0(N1454), 
        .C1(n4306), .Y(n4483) );
  AOI22X1 U4294 ( .A0(N1292), .A1(n4303), .B0(N1369), .B1(n4301), .Y(n4481) );
  AOI222XL U4295 ( .A0(N4377), .A1(n4393), .B0(N4189), .B1(n4394), .C0(N4119), 
        .C1(n3000), .Y(n4479) );
  NAND4BX1 U4296 ( .AN(n4484), .B(n4485), .C(n4486), .D(n4487), .Y(n1432) );
  AOI222XL U4297 ( .A0(N6564), .A1(n3240), .B0(N821), .B1(n3001), .C0(n3243), 
        .C1(N2332), .Y(n4487) );
  NOR3BXL U4298 ( .AN(n4488), .B(n4489), .C(n4490), .Y(n4486) );
  OAI22XL U4299 ( .A0(n4849), .A1(n4381), .B0(n4382), .B1(n4491), .Y(n4490) );
  CLKINVX1 U4300 ( .A(N2418), .Y(n4491) );
  OAI22XL U4301 ( .A0(n3711), .A1(n3248), .B0(n3607), .B1(n3246), .Y(n4489) );
  AOI221XL U4302 ( .A0(N2799), .A1(n3560), .B0(N2864), .B1(n3561), .C0(n4492), 
        .Y(n3607) );
  MXI2X1 U4303 ( .A(N2418), .B(N2332), .S0(n3069), .Y(n3711) );
  AOI222XL U4304 ( .A0(n3208), .A1(n4493), .B0(N501), .B1(n4314), .C0(n3241), 
        .C1(n3758), .Y(n4488) );
  CLKMX2X2 U4305 ( .A(N2418), .B(N2332), .S0(n3381), .Y(n3758) );
  CLKINVX1 U4306 ( .A(n3591), .Y(n4493) );
  AOI221XL U4307 ( .A0(N4990), .A1(n3560), .B0(N5035), .B1(n3561), .C0(n4492), 
        .Y(n3591) );
  NOR2X1 U4308 ( .A(n3623), .B(n4849), .Y(n4492) );
  AOI222XL U4309 ( .A0(N958), .A1(n4308), .B0(N881), .B1(n3291), .C0(N1038), 
        .C1(n3292), .Y(n4485) );
  NAND4X1 U4310 ( .A(n4494), .B(n4495), .C(n4496), .D(n4497), .Y(n4484) );
  AND3X1 U4311 ( .A(n4498), .B(n4499), .C(n4500), .Y(n4497) );
  AOI222XL U4312 ( .A0(N723), .A1(n4304), .B0(N658), .B1(n3013), .C0(N1455), 
        .C1(n4306), .Y(n4500) );
  AOI22X1 U4313 ( .A0(N1293), .A1(n4303), .B0(N1370), .B1(n4301), .Y(n4498) );
  AOI222XL U4314 ( .A0(N4378), .A1(n4393), .B0(N4190), .B1(n4394), .C0(N4120), 
        .C1(n3000), .Y(n4496) );
  NAND4BX1 U4315 ( .AN(n4501), .B(n4502), .C(n4503), .D(n4504), .Y(n1431) );
  AOI222XL U4316 ( .A0(N6565), .A1(n3240), .B0(N822), .B1(n3001), .C0(n3243), 
        .C1(N2333), .Y(n4504) );
  NOR3BXL U4317 ( .AN(n4505), .B(n4506), .C(n4507), .Y(n4503) );
  OAI22XL U4318 ( .A0(n4848), .A1(n4381), .B0(n4382), .B1(n4508), .Y(n4507) );
  CLKINVX1 U4319 ( .A(N2419), .Y(n4508) );
  OAI22XL U4320 ( .A0(n3699), .A1(n3248), .B0(n3617), .B1(n3246), .Y(n4506) );
  AOI221XL U4321 ( .A0(N2800), .A1(n3560), .B0(N2865), .B1(n3561), .C0(n4509), 
        .Y(n3617) );
  AOI222XL U4322 ( .A0(n3208), .A1(n4510), .B0(N502), .B1(n4314), .C0(n3241), 
        .C1(n3746), .Y(n4505) );
  CLKMX2X2 U4323 ( .A(N2419), .B(N2333), .S0(n3381), .Y(n3746) );
  CLKINVX1 U4324 ( .A(n3579), .Y(n4510) );
  AOI221XL U4325 ( .A0(N4991), .A1(n3560), .B0(N5036), .B1(n3561), .C0(n4509), 
        .Y(n3579) );
  NOR2X1 U4326 ( .A(n3623), .B(n4848), .Y(n4509) );
  AOI222XL U4327 ( .A0(N959), .A1(n4308), .B0(N882), .B1(n3291), .C0(N1039), 
        .C1(n3292), .Y(n4502) );
  NAND4X1 U4328 ( .A(n4511), .B(n4512), .C(n4513), .D(n4514), .Y(n4501) );
  AND3X1 U4329 ( .A(n4515), .B(n4516), .C(n4517), .Y(n4514) );
  AOI222XL U4330 ( .A0(N724), .A1(n4304), .B0(N659), .B1(n3013), .C0(N1456), 
        .C1(n4306), .Y(n4517) );
  AOI22X1 U4331 ( .A0(N1294), .A1(n4303), .B0(N1371), .B1(n4301), .Y(n4515) );
  AOI222XL U4332 ( .A0(N4379), .A1(n4393), .B0(N4191), .B1(n4394), .C0(N4121), 
        .C1(n3000), .Y(n4513) );
  NAND4BX1 U4333 ( .AN(n4518), .B(n4519), .C(n4520), .D(n4521), .Y(n1430) );
  AOI222XL U4334 ( .A0(N6566), .A1(n3240), .B0(N823), .B1(n3001), .C0(n3243), 
        .C1(N2334), .Y(n4521) );
  NOR3BXL U4335 ( .AN(n4522), .B(n4523), .C(n4524), .Y(n4520) );
  OAI22XL U4336 ( .A0(n4847), .A1(n4381), .B0(n4382), .B1(n4525), .Y(n4524) );
  CLKINVX1 U4337 ( .A(N2420), .Y(n4525) );
  OAI22XL U4338 ( .A0(n3680), .A1(n3248), .B0(n3635), .B1(n3246), .Y(n4523) );
  AOI221XL U4339 ( .A0(N2801), .A1(n3560), .B0(N2866), .B1(n3561), .C0(n4526), 
        .Y(n3635) );
  AOI222XL U4340 ( .A0(n3208), .A1(n4527), .B0(N503), .B1(n4314), .C0(n3241), 
        .C1(n3727), .Y(n4522) );
  CLKMX2X2 U4341 ( .A(N2420), .B(N2334), .S0(n3381), .Y(n3727) );
  CLKINVX1 U4342 ( .A(n3555), .Y(n4527) );
  AOI221XL U4343 ( .A0(N4992), .A1(n3560), .B0(N5037), .B1(n3561), .C0(n4526), 
        .Y(n3555) );
  NOR2X1 U4344 ( .A(n3623), .B(n4847), .Y(n4526) );
  AOI222XL U4345 ( .A0(N960), .A1(n4308), .B0(N883), .B1(n3291), .C0(N1040), 
        .C1(n3292), .Y(n4519) );
  NAND4X1 U4346 ( .A(n4528), .B(n4529), .C(n4530), .D(n4531), .Y(n4518) );
  AND3X1 U4347 ( .A(n4532), .B(n4533), .C(n4534), .Y(n4531) );
  AOI222XL U4348 ( .A0(N725), .A1(n4304), .B0(N660), .B1(n3013), .C0(N1457), 
        .C1(n4306), .Y(n4534) );
  AOI22X1 U4349 ( .A0(N1295), .A1(n4303), .B0(N1372), .B1(n4301), .Y(n4532) );
  AOI222XL U4350 ( .A0(N4380), .A1(n4393), .B0(N4192), .B1(n4394), .C0(N4122), 
        .C1(n3000), .Y(n4530) );
  NAND4BX1 U4351 ( .AN(n4535), .B(n4536), .C(n4537), .D(n4538), .Y(n1429) );
  AOI222XL U4352 ( .A0(N6567), .A1(n3240), .B0(N824), .B1(n3001), .C0(n3243), 
        .C1(N2335), .Y(n4538) );
  NOR3BXL U4353 ( .AN(n4539), .B(n4540), .C(n4541), .Y(n4537) );
  OAI22XL U4354 ( .A0(n4846), .A1(n4381), .B0(n4382), .B1(n4542), .Y(n4541) );
  CLKINVX1 U4355 ( .A(N2421), .Y(n4542) );
  OAI22XL U4356 ( .A0(n3674), .A1(n3248), .B0(n3639), .B1(n3246), .Y(n4540) );
  AOI221XL U4357 ( .A0(N2802), .A1(n3560), .B0(N2867), .B1(n3561), .C0(n4543), 
        .Y(n3639) );
  MXI2X1 U4358 ( .A(N2421), .B(N2335), .S0(n3069), .Y(n3674) );
  AOI222XL U4359 ( .A0(n3208), .A1(n3548), .B0(N504), .B1(n4314), .C0(n3241), 
        .C1(n3721), .Y(n4539) );
  CLKMX2X2 U4360 ( .A(N2421), .B(N2335), .S0(n3381), .Y(n3721) );
  CLKINVX1 U4361 ( .A(n4544), .Y(n3548) );
  AOI221XL U4362 ( .A0(N4993), .A1(n3560), .B0(N5038), .B1(n3561), .C0(n4543), 
        .Y(n4544) );
  NOR2X1 U4363 ( .A(n3623), .B(n4846), .Y(n4543) );
  AOI222XL U4364 ( .A0(N961), .A1(n4308), .B0(N884), .B1(n3291), .C0(N1041), 
        .C1(n3292), .Y(n4536) );
  NAND4X1 U4365 ( .A(n4545), .B(n4546), .C(n4547), .D(n4548), .Y(n4535) );
  AND3X1 U4366 ( .A(n4549), .B(n4550), .C(n4551), .Y(n4548) );
  AOI222XL U4367 ( .A0(N726), .A1(n4304), .B0(N661), .B1(n3013), .C0(N1458), 
        .C1(n4306), .Y(n4551) );
  AOI22X1 U4368 ( .A0(N1296), .A1(n4303), .B0(N1373), .B1(n4301), .Y(n4549) );
  AOI222XL U4369 ( .A0(N4381), .A1(n4393), .B0(N4193), .B1(n4394), .C0(N4123), 
        .C1(n3000), .Y(n4547) );
  NAND4BX1 U4370 ( .AN(n4552), .B(n4553), .C(n4554), .D(n4555), .Y(n1428) );
  AOI222XL U4371 ( .A0(N6568), .A1(n3240), .B0(N825), .B1(n3001), .C0(n3243), 
        .C1(N2336), .Y(n4555) );
  NOR3BXL U4372 ( .AN(n4556), .B(n4557), .C(n4558), .Y(n4554) );
  OAI22XL U4373 ( .A0(n4845), .A1(n4381), .B0(n4382), .B1(n4559), .Y(n4558) );
  CLKINVX1 U4374 ( .A(N2422), .Y(n4559) );
  OAI22XL U4375 ( .A0(n3676), .A1(n3248), .B0(n3637), .B1(n3246), .Y(n4557) );
  AOI221XL U4376 ( .A0(N2803), .A1(n3560), .B0(N2868), .B1(n3561), .C0(n4560), 
        .Y(n3637) );
  MXI2X1 U4377 ( .A(N2422), .B(N2336), .S0(n3069), .Y(n3676) );
  AOI222XL U4378 ( .A0(n3208), .A1(n3550), .B0(N505), .B1(n4314), .C0(n3241), 
        .C1(n3723), .Y(n4556) );
  CLKMX2X2 U4379 ( .A(N2422), .B(N2336), .S0(n3381), .Y(n3723) );
  CLKINVX1 U4380 ( .A(n4561), .Y(n3550) );
  AOI221XL U4381 ( .A0(N4994), .A1(n3560), .B0(N5039), .B1(n3561), .C0(n4560), 
        .Y(n4561) );
  NOR2X1 U4382 ( .A(n3623), .B(n4845), .Y(n4560) );
  AOI222XL U4383 ( .A0(N962), .A1(n4308), .B0(N885), .B1(n3291), .C0(N1042), 
        .C1(n3292), .Y(n4553) );
  NAND4X1 U4384 ( .A(n4562), .B(n4563), .C(n4564), .D(n4565), .Y(n4552) );
  AND3X1 U4385 ( .A(n4566), .B(n4567), .C(n4568), .Y(n4565) );
  AOI222XL U4386 ( .A0(N727), .A1(n4304), .B0(N662), .B1(n3013), .C0(N1459), 
        .C1(n4306), .Y(n4568) );
  AOI22X1 U4387 ( .A0(N1297), .A1(n4303), .B0(N1374), .B1(n4301), .Y(n4566) );
  AOI222XL U4388 ( .A0(N4382), .A1(n4393), .B0(N4194), .B1(n4394), .C0(N4124), 
        .C1(n3000), .Y(n4564) );
  NAND4BX1 U4389 ( .AN(n4569), .B(n4570), .C(n4571), .D(n4572), .Y(n1427) );
  AOI222XL U4390 ( .A0(N6569), .A1(n3240), .B0(n3241), .B1(n3722), .C0(n3208), 
        .C1(n3549), .Y(n4572) );
  CLKINVX1 U4391 ( .A(n4573), .Y(n3549) );
  AOI221XL U4392 ( .A0(N4995), .A1(n3560), .B0(N5040), .B1(n3561), .C0(n4574), 
        .Y(n4573) );
  CLKMX2X2 U4393 ( .A(N2423), .B(N2337), .S0(n3381), .Y(n3722) );
  NOR3BXL U4394 ( .AN(n4575), .B(n4576), .C(n4577), .Y(n4571) );
  OAI22XL U4395 ( .A0(n4844), .A1(n4381), .B0(n4382), .B1(n4578), .Y(n4577) );
  CLKINVX1 U4396 ( .A(N2423), .Y(n4578) );
  OAI22XL U4397 ( .A0(n3675), .A1(n3248), .B0(n3638), .B1(n3246), .Y(n4576) );
  AOI221XL U4398 ( .A0(N2804), .A1(n3560), .B0(N2869), .B1(n3561), .C0(n4574), 
        .Y(n3638) );
  NOR2X1 U4399 ( .A(n3623), .B(n4844), .Y(n4574) );
  MXI2X1 U4400 ( .A(N2423), .B(N2337), .S0(n3069), .Y(n3675) );
  AOI222XL U4401 ( .A0(N1043), .A1(n3292), .B0(N506), .B1(n4314), .C0(N886), 
        .C1(n3291), .Y(n4575) );
  AOI222XL U4402 ( .A0(n3243), .A1(N2337), .B0(N963), .B1(n4308), .C0(N826), 
        .C1(n3001), .Y(n4570) );
  NAND4X1 U4403 ( .A(n4581), .B(n4582), .C(n4583), .D(n4584), .Y(n4569) );
  AND3X1 U4404 ( .A(n4585), .B(n4586), .C(n4587), .Y(n4584) );
  AOI222XL U4405 ( .A0(N728), .A1(n4304), .B0(N663), .B1(n3013), .C0(N1460), 
        .C1(n4306), .Y(n4587) );
  AOI22X1 U4406 ( .A0(N527), .A1(n4300), .B0(N567), .B1(n4302), .Y(n4586) );
  AOI22X1 U4407 ( .A0(N1298), .A1(n4303), .B0(N1375), .B1(n4301), .Y(n4585) );
  AOI222XL U4408 ( .A0(N4383), .A1(n4393), .B0(N4195), .B1(n4394), .C0(N4125), 
        .C1(n3000), .Y(n4583) );
  NAND3X1 U4409 ( .A(n4588), .B(n4589), .C(n4590), .Y(n1426) );
  NOR4X1 U4410 ( .A(n4591), .B(n4592), .C(n4593), .D(n4594), .Y(n4590) );
  AO22X1 U4411 ( .A0(N1026), .A1(n3292), .B0(N869), .B1(n3291), .Y(n4594) );
  NAND2X1 U4412 ( .A(n3468), .B(n3561), .Y(n3259) );
  NAND2X1 U4413 ( .A(n3469), .B(n3561), .Y(n3258) );
  OAI2BB2XL U4414 ( .B0(n3700), .B1(n3248), .A0N(n4286), .A1N(N489), .Y(n4593)
         );
  CLKINVX1 U4415 ( .A(n3293), .Y(n4286) );
  NAND2X1 U4416 ( .A(n3371), .B(n3255), .Y(n3293) );
  CLKINVX1 U4417 ( .A(n3442), .Y(n3255) );
  NAND2X1 U4418 ( .A(n2016), .B(n3372), .Y(n3442) );
  NAND2X1 U4419 ( .A(n3343), .B(n3531), .Y(n3328) );
  MXI2X1 U4420 ( .A(N3734), .B(N2320), .S0(n3069), .Y(n3700) );
  OAI2BB2XL U4421 ( .B0(n3618), .B1(n3246), .A0N(N3734), .A1N(n3195), .Y(n4592) );
  NAND2X1 U4422 ( .A(n3422), .B(n2979), .Y(n3331) );
  CLKINVX1 U4423 ( .A(n3417), .Y(n3336) );
  NAND2X1 U4424 ( .A(n3449), .B(n3531), .Y(n3417) );
  AOI221XL U4425 ( .A0(N2787), .A1(n3560), .B0(N2852), .B1(n3561), .C0(n4595), 
        .Y(n3618) );
  OAI222XL U4426 ( .A0(n3284), .A1(n4596), .B0(n4874), .B1(n3199), .C0(n3286), 
        .C1(n4597), .Y(n4591) );
  CLKINVX1 U4427 ( .A(N946), .Y(n4597) );
  NAND2X1 U4428 ( .A(n3234), .B(n3371), .Y(n3286) );
  CLKINVX1 U4429 ( .A(N809), .Y(n4596) );
  NAND2X1 U4430 ( .A(n3210), .B(n3234), .Y(n3284) );
  CLKINVX1 U4431 ( .A(n4260), .Y(n3234) );
  NAND2X1 U4432 ( .A(n3469), .B(n3560), .Y(n4260) );
  CLKINVX1 U4433 ( .A(n4598), .Y(n3469) );
  NOR4X1 U4434 ( .A(n4599), .B(n4600), .C(n4601), .D(n4602), .Y(n4589) );
  NOR2X1 U4435 ( .A(n3747), .B(n3297), .Y(n4602) );
  NAND2X1 U4436 ( .A(n3343), .B(n3410), .Y(n3297) );
  MXI2X1 U4437 ( .A(N2320), .B(N3734), .S0(n3069), .Y(n3747) );
  AOI21X1 U4438 ( .A0(n4603), .A1(n4604), .B0(n3244), .Y(n4601) );
  AOI222XL U4439 ( .A0(N646), .A1(n3237), .B0(N510), .B1(n3254), .C0(N550), 
        .C1(n3257), .Y(n4604) );
  NOR2BX1 U4440 ( .AN(n4236), .B(n3946), .Y(n3257) );
  NOR2BX1 U4441 ( .AN(n4236), .B(n3950), .Y(n3254) );
  NOR2X1 U4442 ( .A(n3451), .B(n2016), .Y(n4236) );
  AOI22X1 U4443 ( .A0(N711), .A1(n3238), .B0(N809), .B1(n3239), .Y(n4603) );
  OAI2BB2XL U4444 ( .B0(n4842), .B1(n3290), .A0N(N2320), .A1N(n3243), .Y(n4600) );
  NAND2X1 U4445 ( .A(n3422), .B(n2016), .Y(n3665) );
  AOI221XL U4446 ( .A0(n3371), .A1(n3256), .B0(n3210), .B1(n3233), .C0(n3206), 
        .Y(n4607) );
  AOI2BB2X1 U4447 ( .B0(n3406), .B1(state[0]), .A0N(n4264), .A1N(n4608), .Y(
        n3206) );
  NOR2X1 U4448 ( .A(n2963), .B(n2957), .Y(n4264) );
  NAND2X1 U4449 ( .A(n3623), .B(n4243), .Y(n3233) );
  OAI211X1 U4450 ( .A0(n3623), .A1(n4598), .B0(n4243), .C0(n4609), .Y(n3256)
         );
  AOI2BB1X1 U4451 ( .A0N(n3623), .A1N(n3383), .B0(n4242), .Y(n4609) );
  CLKINVX1 U4452 ( .A(n4210), .Y(n4242) );
  NAND2X1 U4453 ( .A(n3449), .B(n4202), .Y(n4210) );
  NAND2X1 U4454 ( .A(n3343), .B(n3381), .Y(n4598) );
  AOI221XL U4455 ( .A0(n3319), .A1(n4610), .B0(n3205), .B1(n4611), .C0(n3207), 
        .Y(n4606) );
  OAI211X1 U4456 ( .A0(n3201), .A1(n3527), .B0(n3407), .C0(n4211), .Y(n3207)
         );
  NAND2BX1 U4457 ( .AN(n4217), .B(n3340), .Y(n4211) );
  NAND2X1 U4458 ( .A(n4001), .B(n4605), .Y(n3407) );
  CLKINVX1 U4459 ( .A(n4610), .Y(n3201) );
  NAND2X1 U4460 ( .A(n3531), .B(n4243), .Y(n4610) );
  NAND2X1 U4461 ( .A(n3375), .B(n3415), .Y(n4243) );
  CLKINVX1 U4462 ( .A(n3396), .Y(n3375) );
  NAND2X1 U4463 ( .A(n3379), .B(n3451), .Y(n3396) );
  AOI21X1 U4464 ( .A0(n4612), .A1(n4613), .B0(n3376), .Y(n4599) );
  NAND2X1 U4465 ( .A(n4001), .B(n3531), .Y(n3463) );
  AOI222XL U4466 ( .A0(N1358), .A1(n3237), .B0(N1281), .B1(n3235), .C0(N489), 
        .C1(n3236), .Y(n4613) );
  CLKINVX1 U4467 ( .A(n4580), .Y(n3236) );
  NAND2X1 U4468 ( .A(n3560), .B(n3372), .Y(n4580) );
  AOI22X1 U4469 ( .A0(N1443), .A1(n3238), .B0(N946), .B1(n3239), .Y(n4612) );
  CLKINVX1 U4470 ( .A(n3270), .Y(n3239) );
  CLKINVX1 U4471 ( .A(n3383), .Y(n3468) );
  AOI211X1 U4472 ( .A0(N6552), .A1(n3240), .B0(n4614), .C0(n4615), .Y(n4588)
         );
  MXI2X1 U4473 ( .A(n4282), .B(n4616), .S0(n4787), .Y(n4615) );
  OR2X1 U4474 ( .A(n3200), .B(n4788), .Y(n4616) );
  OA21XL U4475 ( .A0(n3200), .A1(n2981), .B0(n3289), .Y(n4282) );
  NAND2X1 U4476 ( .A(n3356), .B(n3423), .Y(n3289) );
  CLKINVX1 U4477 ( .A(n3365), .Y(n3423) );
  NAND2X1 U4478 ( .A(n3205), .B(n4251), .Y(n3200) );
  CLKINVX1 U4479 ( .A(n4611), .Y(n4251) );
  NAND2X1 U4480 ( .A(n3787), .B(n3818), .Y(n4611) );
  NOR2X1 U4481 ( .A(n3365), .B(n3356), .Y(n3205) );
  CLKINVX1 U4482 ( .A(n3438), .Y(n3356) );
  NAND2X1 U4483 ( .A(n3818), .B(n4223), .Y(n3438) );
  NOR2X1 U4484 ( .A(N6483), .B(n1424), .Y(n4223) );
  OAI2BB2XL U4485 ( .B0(n3295), .B1(n3580), .A0N(n3212), .A1N(n4617), .Y(n4614) );
  NAND4X1 U4486 ( .A(n4618), .B(n4619), .C(n4620), .D(n4621), .Y(n4617) );
  AOI222XL U4487 ( .A0(N3754), .A1(n3218), .B0(n3219), .B1(IM_A[2]), .C0(N3619), .C1(n3220), .Y(n4621) );
  OAI21XL U4488 ( .A0(n3766), .A1(n4209), .B0(n4257), .Y(n4579) );
  CLKINVX1 U4489 ( .A(n4023), .Y(n4209) );
  AOI22X1 U4490 ( .A0(N3734), .A1(n3221), .B0(N3734), .B1(n3222), .Y(n4620) );
  NAND3X1 U4491 ( .A(\gt_332/n15 ), .B(n3305), .C(n4857), .Y(n3990) );
  NAND3X1 U4492 ( .A(n4857), .B(\gt_332/n15 ), .C(n4855), .Y(n4004) );
  CLKINVX1 U4493 ( .A(n3761), .Y(n3766) );
  NAND2X1 U4494 ( .A(n3595), .B(n3425), .Y(n3712) );
  AND4X1 U4495 ( .A(count[4]), .B(n3424), .C(count[3]), .D(n4623), .Y(n3595)
         );
  NOR2X1 U4496 ( .A(n4874), .B(n4875), .Y(n4623) );
  CLKINVX1 U4497 ( .A(n3436), .Y(n3212) );
  AOI221XL U4498 ( .A0(N4978), .A1(n3560), .B0(N5023), .B1(n3561), .C0(n4595), 
        .Y(n3580) );
  NOR2X1 U4499 ( .A(n3623), .B(n4842), .Y(n4595) );
  NOR2X1 U4500 ( .A(n3560), .B(n3561), .Y(n4202) );
  NAND2X1 U4501 ( .A(n4856), .B(n4857), .Y(n4257) );
  NAND2X1 U4502 ( .A(n3449), .B(n3410), .Y(n3295) );
  NOR4X1 U4503 ( .A(pic_size[6]), .B(pic_size[5]), .C(pic_size[4]), .D(
        pic_size[3]), .Y(n4624) );
  CLKINVX1 U4504 ( .A(n3527), .Y(n3360) );
  NAND2X1 U4505 ( .A(n3367), .B(n3478), .Y(n3527) );
  OAI21XL U4506 ( .A0(n3787), .A1(n4874), .B0(n4258), .Y(n4625) );
  CLKINVX1 U4507 ( .A(reset), .Y(n1425) );
  OAI22XL U4508 ( .A0(n4626), .A1(n4627), .B0(n4628), .B1(n4629), .Y(min_n[6])
         );
  CLKINVX1 U4509 ( .A(N6789), .Y(n4627) );
  OAI222XL U4510 ( .A0(n4628), .A1(n4630), .B0(n4864), .B1(n4631), .C0(n4632), 
        .C1(n4626), .Y(min_n[5]) );
  CLKINVX1 U4511 ( .A(N6788), .Y(n4632) );
  OAI222XL U4512 ( .A0(n4866), .A1(n4631), .B0(n3814), .B1(n4633), .C0(n4634), 
        .C1(n4626), .Y(min_n[4]) );
  CLKINVX1 U4513 ( .A(N6787), .Y(n4634) );
  CLKINVX1 U4514 ( .A(IM_Q[12]), .Y(n3814) );
  OAI222XL U4515 ( .A0(n4868), .A1(n4631), .B0(n3815), .B1(n4633), .C0(n4635), 
        .C1(n4626), .Y(min_n[3]) );
  CLKINVX1 U4516 ( .A(N6786), .Y(n4635) );
  CLKINVX1 U4517 ( .A(IM_Q[11]), .Y(n3815) );
  OAI222XL U4518 ( .A0(n4867), .A1(n4631), .B0(n3816), .B1(n4633), .C0(n4636), 
        .C1(n4626), .Y(min_n[2]) );
  NAND2X1 U4519 ( .A(n4637), .B(n4638), .Y(n4633) );
  CLKINVX1 U4520 ( .A(IM_Q[10]), .Y(n3816) );
  NAND2X1 U4521 ( .A(n4639), .B(n4638), .Y(n4631) );
  OAI22XL U4522 ( .A0(n4626), .A1(n4640), .B0(n4628), .B1(n4641), .Y(min_n[1])
         );
  CLKINVX1 U4523 ( .A(N6784), .Y(n4640) );
  OAI22XL U4524 ( .A0(n4626), .A1(n4642), .B0(n4628), .B1(n4643), .Y(min_n[0])
         );
  CLKINVX1 U4525 ( .A(n4638), .Y(n4628) );
  CLKINVX1 U4526 ( .A(N6783), .Y(n4642) );
  OAI22XL U4527 ( .A0(n4646), .A1(n4647), .B0(n4648), .B1(n4649), .Y(hour_n[6]) );
  CLKINVX1 U4528 ( .A(n4650), .Y(n4649) );
  CLKINVX1 U4529 ( .A(N6810), .Y(n4647) );
  OAI22XL U4530 ( .A0(n4646), .A1(n4651), .B0(n4648), .B1(n4652), .Y(hour_n[5]) );
  CLKINVX1 U4531 ( .A(n4653), .Y(n4652) );
  CLKINVX1 U4532 ( .A(N6809), .Y(n4651) );
  OAI22XL U4533 ( .A0(n4654), .A1(n4646), .B0(n4648), .B1(n4655), .Y(hour_n[4]) );
  OA22X1 U4534 ( .A0(n3996), .A1(n4656), .B0(n4657), .B1(n4861), .Y(n4655) );
  CLKINVX1 U4535 ( .A(IM_Q[20]), .Y(n3996) );
  CLKINVX1 U4536 ( .A(N6808), .Y(n4654) );
  OAI22XL U4537 ( .A0(n4658), .A1(n4646), .B0(n4648), .B1(n4659), .Y(hour_n[3]) );
  OA21XL U4538 ( .A0(n3806), .A1(n4656), .B0(n4660), .Y(n4659) );
  CLKINVX1 U4539 ( .A(N6807), .Y(n4658) );
  OAI22XL U4540 ( .A0(n4646), .A1(n4661), .B0(n4648), .B1(n4662), .Y(hour_n[2]) );
  CLKINVX1 U4541 ( .A(n4663), .Y(n4662) );
  CLKINVX1 U4542 ( .A(N6806), .Y(n4661) );
  OAI22XL U4543 ( .A0(n4646), .A1(n4664), .B0(n4648), .B1(n4665), .Y(hour_n[1]) );
  CLKINVX1 U4544 ( .A(n4666), .Y(n4665) );
  CLKINVX1 U4545 ( .A(N6805), .Y(n4664) );
  OAI22XL U4546 ( .A0(n4646), .A1(n4667), .B0(n4648), .B1(n4668), .Y(hour_n[0]) );
  MXI2X1 U4547 ( .A(n4670), .B(n4671), .S0(n4645), .Y(n4669) );
  CLKINVX1 U4548 ( .A(n3783), .Y(n4644) );
  NAND4X1 U4549 ( .A(N6773), .B(N6772), .C(N6774), .D(n4674), .Y(n3783) );
  NOR4X1 U4550 ( .A(N6775), .B(N6770), .C(N6769), .D(n3777), .Y(n4674) );
  CLKINVX1 U4551 ( .A(N6771), .Y(n3777) );
  NAND4X1 U4552 ( .A(N6787), .B(N6786), .C(N6788), .D(n4675), .Y(n4673) );
  NOR4X1 U4553 ( .A(N6789), .B(N6784), .C(N6783), .D(n4636), .Y(n4675) );
  CLKINVX1 U4554 ( .A(N6785), .Y(n4636) );
  NAND4X1 U4555 ( .A(n4641), .B(n4643), .C(n4629), .D(n4676), .Y(n4672) );
  AOI222XL U4556 ( .A0(n3982), .A1(n4656), .B0(n4864), .B1(n4630), .C0(n4657), 
        .C1(n4677), .Y(n4676) );
  NAND4BX1 U4557 ( .AN(n4630), .B(IM_Q[10]), .C(IM_Q[11]), .D(IM_Q[12]), .Y(
        n4677) );
  NAND2X1 U4558 ( .A(n4637), .B(IM_Q[13]), .Y(n4630) );
  CLKINVX1 U4559 ( .A(n4656), .Y(n4637) );
  NAND3X1 U4560 ( .A(n3979), .B(min[4]), .C(n3980), .Y(n3982) );
  CLKINVX1 U4561 ( .A(n4868), .Y(n3980) );
  CLKINVX1 U4562 ( .A(n4867), .Y(n3979) );
  OA22X1 U4563 ( .A0(n3812), .A1(n4656), .B0(n4865), .B1(n4657), .Y(n4629) );
  CLKINVX1 U4564 ( .A(IM_Q[14]), .Y(n3812) );
  AOI2BB2X1 U4565 ( .B0(N6150), .B1(n4639), .A0N(n3470), .A1N(n4656), .Y(n4641) );
  NAND4X1 U4566 ( .A(N6807), .B(n4667), .C(N6808), .D(n4678), .Y(n4671) );
  NOR4X1 U4567 ( .A(N6810), .B(N6809), .C(N6806), .D(N6805), .Y(n4678) );
  CLKINVX1 U4568 ( .A(N6804), .Y(n4667) );
  NAND4X1 U4569 ( .A(n4679), .B(n4680), .C(n4681), .D(n4682), .Y(n4670) );
  NOR4X1 U4570 ( .A(n4666), .B(n4663), .C(n4653), .D(n4650), .Y(n4682) );
  OAI22XL U4571 ( .A0(n4860), .A1(n4657), .B0(n3994), .B1(n4656), .Y(n4650) );
  CLKINVX1 U4572 ( .A(IM_Q[22]), .Y(n3994) );
  OAI22XL U4573 ( .A0(n4859), .A1(n4657), .B0(n3995), .B1(n4656), .Y(n4653) );
  CLKINVX1 U4574 ( .A(IM_Q[21]), .Y(n3995) );
  OAI22XL U4575 ( .A0(n4863), .A1(n4657), .B0(n3808), .B1(n4656), .Y(n4663) );
  CLKINVX1 U4576 ( .A(IM_Q[18]), .Y(n3808) );
  OAI22XL U4577 ( .A0(n4858), .A1(n4657), .B0(n3809), .B1(n4656), .Y(n4666) );
  CLKINVX1 U4578 ( .A(IM_Q[17]), .Y(n3809) );
  OA21XL U4579 ( .A0(IM_Q[20]), .A1(n4639), .B0(n4668), .Y(n4681) );
  OA22X1 U4580 ( .A0(n3810), .A1(n4656), .B0(n4809), .B1(n4657), .Y(n4668) );
  CLKINVX1 U4581 ( .A(IM_Q[16]), .Y(n3810) );
  OAI21XL U4582 ( .A0(n3806), .A1(n4656), .B0(n4660), .Y(n4680) );
  NAND2BX1 U4583 ( .AN(n4862), .B(n4639), .Y(n4660) );
  OAI211X1 U4584 ( .A0(n3781), .A1(n3199), .B0(n3805), .C0(n4683), .Y(n4639)
         );
  NOR2X1 U4585 ( .A(n3367), .B(n3370), .Y(n4683) );
  CLKINVX1 U4586 ( .A(n3325), .Y(n3370) );
  NAND2X1 U4587 ( .A(state[2]), .B(state[1]), .Y(n3325) );
  NAND2X1 U4588 ( .A(n4263), .B(state[0]), .Y(n3798) );
  AND4X1 U4589 ( .A(n3457), .B(n3365), .C(n3406), .D(n4684), .Y(n3805) );
  NOR2X1 U4590 ( .A(n3357), .B(n4001), .Y(n4684) );
  CLKINVX1 U4591 ( .A(n3458), .Y(n4001) );
  NAND2X1 U4592 ( .A(n4263), .B(n2973), .Y(n3458) );
  NOR2X1 U4593 ( .A(n2957), .B(state[2]), .Y(n4263) );
  NAND3X1 U4594 ( .A(state[2]), .B(state[1]), .C(state[0]), .Y(n3406) );
  NAND3X1 U4595 ( .A(n2957), .B(n2963), .C(state[0]), .Y(n3365) );
  NAND2X1 U4596 ( .A(n4608), .B(state[0]), .Y(n3457) );
  NOR2X1 U4597 ( .A(n2963), .B(state[1]), .Y(n4608) );
  NAND2X1 U4598 ( .A(n4861), .B(n4656), .Y(n4679) );
  NAND3X1 U4599 ( .A(n2957), .B(n2963), .C(n2973), .Y(n3199) );
  AND2X1 U4600 ( .A(n4225), .B(n3818), .Y(n3781) );
  NOR2X1 U4601 ( .A(N6484), .B(n3788), .Y(n3818) );
  NAND2X1 U4602 ( .A(n4873), .B(n4258), .Y(n3788) );
  NOR4X1 U4603 ( .A(n3425), .B(n3426), .C(n3424), .D(count[4]), .Y(n4258) );
  CLKINVX1 U4604 ( .A(n4872), .Y(n3424) );
  CLKINVX1 U4605 ( .A(n4871), .Y(n3426) );
  CLKINVX1 U4606 ( .A(n4870), .Y(n3425) );
  NOR2X1 U4607 ( .A(n3188), .B(n4875), .Y(n4225) );
  CLKINVX1 U4608 ( .A(n1424), .Y(n3188) );
  AND2X1 U4609 ( .A(N6754), .B(n3187), .Y(cycle_n[9]) );
  AND2X1 U4610 ( .A(N6753), .B(n3187), .Y(cycle_n[8]) );
  AND2X1 U4611 ( .A(N6752), .B(n3187), .Y(cycle_n[7]) );
  AND2X1 U4612 ( .A(N6751), .B(n3187), .Y(cycle_n[6]) );
  AND2X1 U4613 ( .A(N6750), .B(n3187), .Y(cycle_n[5]) );
  AND2X1 U4614 ( .A(N6749), .B(n3187), .Y(cycle_n[4]) );
  AND2X1 U4615 ( .A(N6748), .B(n3187), .Y(cycle_n[3]) );
  AND2X1 U4616 ( .A(N6747), .B(n3187), .Y(cycle_n[2]) );
  AND2X1 U4617 ( .A(N6746), .B(n3187), .Y(cycle_n[1]) );
  AND2X1 U4618 ( .A(N6764), .B(n3187), .Y(cycle_n[19]) );
  AND2X1 U4619 ( .A(N6763), .B(n3187), .Y(cycle_n[18]) );
  AND2X1 U4620 ( .A(N6762), .B(n3187), .Y(cycle_n[17]) );
  AND2X1 U4621 ( .A(N6761), .B(n3187), .Y(cycle_n[16]) );
  AND2X1 U4622 ( .A(N6760), .B(n3187), .Y(cycle_n[15]) );
  AND2X1 U4623 ( .A(N6759), .B(n3187), .Y(cycle_n[14]) );
  AND2X1 U4624 ( .A(N6758), .B(n3187), .Y(cycle_n[13]) );
  AND2X1 U4625 ( .A(N6757), .B(n3187), .Y(cycle_n[12]) );
  AND2X1 U4626 ( .A(N6756), .B(n3187), .Y(cycle_n[11]) );
  AND2X1 U4627 ( .A(N6755), .B(n3187), .Y(cycle_n[10]) );
  AND2X1 U4628 ( .A(N6745), .B(n3187), .Y(cycle_n[0]) );
  NOR4X1 U4629 ( .A(n4689), .B(n4690), .C(n4691), .D(n4692), .Y(n4688) );
  NOR3X1 U4630 ( .A(n4699), .B(n4694), .C(n4697), .Y(n4687) );
  NOR4X1 U4631 ( .A(n4700), .B(n4705), .C(n4706), .D(n4744), .Y(n4686) );
  NOR3X1 U4632 ( .A(n3804), .B(n4745), .C(n3799), .Y(n4685) );
  NAND4X1 U4633 ( .A(n4701), .B(n4702), .C(n4703), .D(n4704), .Y(n3799) );
  NAND4X1 U4634 ( .A(n4693), .B(n4695), .C(n4696), .D(n4698), .Y(n3804) );
endmodule

